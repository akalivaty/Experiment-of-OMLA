//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n590, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT65), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(KEYINPUT65), .B1(G567), .B2(new_n453), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n462), .A2(new_n464), .A3(new_n468), .A4(new_n465), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(G2104), .B2(new_n468), .ZN(new_n474));
  NOR3_X1   g049(.A1(new_n461), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(G101), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G101), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n469), .A2(new_n472), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n463), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(new_n465), .A3(G125), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(KEYINPUT66), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n486), .B(new_n468), .C1(new_n482), .C2(new_n483), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  INV_X1    g065(.A(G100), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n491), .A2(new_n468), .A3(KEYINPUT71), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT71), .B1(new_n491), .B2(new_n468), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G112), .B2(new_n468), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G124), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n462), .A2(new_n464), .A3(G2105), .A4(new_n465), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n470), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(G136), .B2(new_n498), .ZN(G162));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  AND4_X1   g077(.A1(G2105), .A2(new_n462), .A3(new_n464), .A4(new_n465), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G126), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n462), .A2(new_n464), .A3(new_n506), .A4(new_n465), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n481), .A2(new_n465), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n505), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n504), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n507), .A2(KEYINPUT4), .B1(new_n509), .B2(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(new_n500), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(G114), .B2(new_n468), .ZN(new_n517));
  INV_X1    g092(.A(G126), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n496), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT72), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(new_n527), .B1(new_n524), .B2(G543), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n529), .A2(G543), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(G88), .B1(G50), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(G62), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n528), .A2(new_n529), .ZN(new_n540));
  INV_X1    g115(.A(G88), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n529), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G50), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n533), .B2(new_n534), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n539), .A2(new_n548), .ZN(G303));
  INV_X1    g124(.A(G303), .ZN(G166));
  NAND2_X1  g125(.A1(new_n531), .A2(G51), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n552));
  NAND3_X1  g127(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n530), .A2(G89), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(G168));
  AOI22_X1  g132(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n545), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  INV_X1    g135(.A(G52), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n540), .A2(new_n560), .B1(new_n542), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(G171));
  AOI22_X1  g138(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n545), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n530), .A2(G81), .B1(G43), .B2(new_n531), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT75), .Z(G176));
  XOR2_X1   g146(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n572));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  XOR2_X1   g150(.A(KEYINPUT78), .B(G65), .Z(new_n576));
  AOI22_X1  g151(.A1(new_n528), .A2(new_n576), .B1(G78), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n545), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT79), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n531), .A2(G53), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(G91), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n540), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n530), .A2(KEYINPUT77), .A3(G91), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n579), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G171), .ZN(G301));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(G168), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n555), .A2(new_n556), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT80), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(G286));
  OAI21_X1  g169(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n531), .A2(G49), .ZN(new_n596));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n540), .ZN(G288));
  AOI22_X1  g173(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n545), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n600), .A2(new_n601), .B1(G48), .B2(new_n531), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT81), .B1(new_n599), .B2(new_n545), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n530), .A2(G86), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(G305));
  AOI22_X1  g183(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n545), .ZN(new_n610));
  INV_X1    g185(.A(G85), .ZN(new_n611));
  INV_X1    g186(.A(G47), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n540), .A2(new_n611), .B1(new_n542), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n530), .A2(G92), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n528), .A2(G66), .ZN(new_n620));
  INV_X1    g195(.A(G79), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n526), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(G54), .B2(new_n531), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n616), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n616), .B1(new_n625), .B2(G868), .ZN(G321));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NOR2_X1   g203(.A1(G286), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n579), .A2(new_n587), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n629), .B1(new_n631), .B2(new_n628), .ZN(G297));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n628), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n625), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND3_X1  g210(.A1(new_n625), .A2(KEYINPUT84), .A3(new_n634), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n624), .B2(G559), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  MUX2_X1   g214(.A(new_n567), .B(new_n639), .S(G868), .Z(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g216(.A(new_n509), .B1(new_n475), .B2(new_n474), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n647));
  INV_X1    g222(.A(G111), .ZN(new_n648));
  AOI22_X1  g223(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(G2105), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n647), .B2(new_n646), .ZN(new_n650));
  INV_X1    g225(.A(G123), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n496), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(G135), .B2(new_n498), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2096), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n645), .A2(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2451), .B(G2454), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n663), .B(new_n666), .Z(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n663), .A2(new_n666), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n663), .A2(new_n666), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n674), .B2(new_n668), .ZN(new_n675));
  AOI211_X1 g250(.A(KEYINPUT87), .B(new_n669), .C1(new_n672), .C2(new_n673), .ZN(new_n676));
  OAI211_X1 g251(.A(G14), .B(new_n670), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(G401));
  XNOR2_X1  g253(.A(KEYINPUT91), .B(G2100), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2084), .B(G2090), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(KEYINPUT17), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n681), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n682), .A2(new_n681), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n687), .B(new_n691), .C1(new_n685), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G2096), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(G2096), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n680), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(new_n694), .A3(new_n679), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(G227));
  XNOR2_X1  g275(.A(G1956), .B(G2474), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT92), .ZN(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1971), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT19), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n706), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n709), .A2(new_n702), .A3(new_n703), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT20), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(KEYINPUT20), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n708), .B1(new_n706), .B2(new_n704), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1991), .B(G1996), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(G1981), .B(G1986), .ZN(new_n720));
  INV_X1    g295(.A(new_n714), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n713), .A2(new_n721), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n722), .A2(new_n723), .A3(new_n717), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n720), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n715), .A2(new_n718), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n724), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n729), .ZN(G229));
  NAND2_X1  g305(.A1(G168), .A2(G16), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(KEYINPUT99), .C1(G16), .C2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(KEYINPUT99), .B2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G1966), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT100), .Z(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  NAND2_X1  g311(.A1(G164), .A2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G27), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G32), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n503), .A2(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(G105), .B1(new_n474), .B2(new_n475), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n498), .A2(G141), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n741), .B1(new_n749), .B2(new_n740), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT97), .Z(new_n751));
  OAI221_X1 g326(.A(new_n735), .B1(new_n736), .B2(new_n738), .C1(new_n739), .C2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n740), .B1(KEYINPUT24), .B2(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n489), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n752), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n753), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n740), .A2(G33), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  AOI22_X1  g337(.A1(new_n509), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n468), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G139), .B2(new_n498), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n760), .B1(new_n765), .B2(new_n740), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2072), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n759), .B(new_n767), .C1(new_n739), .C2(new_n751), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n733), .A2(G1966), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G19), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n568), .B2(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n653), .A2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT30), .B(G28), .ZN(new_n776));
  OR2_X1    g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n776), .A2(new_n740), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n774), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n773), .A2(G1341), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n771), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n738), .A2(new_n736), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n625), .B2(G16), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n740), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  INV_X1    g365(.A(G128), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n468), .A2(G116), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n496), .A2(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n498), .B2(G140), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n790), .B1(new_n795), .B2(new_n740), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G16), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n799), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT101), .B(G1961), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n788), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G29), .A2(G35), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G162), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n799), .A2(G20), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT23), .Z(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G299), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n784), .A2(new_n804), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n758), .A2(new_n770), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n799), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n799), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(G1971), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(G1971), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n799), .A2(G23), .ZN(new_n820));
  INV_X1    g395(.A(G288), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n799), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT33), .B(G1976), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n818), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n799), .A2(G6), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n604), .A2(new_n607), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n799), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT32), .B(G1981), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT94), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n825), .A2(new_n831), .A3(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n799), .A2(G24), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n614), .B2(new_n799), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G1986), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n740), .A2(G25), .ZN(new_n836));
  INV_X1    g411(.A(G119), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n468), .A2(G107), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n496), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n498), .B2(G131), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n836), .B1(new_n841), .B2(new_n740), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  XOR2_X1   g418(.A(new_n842), .B(new_n843), .Z(new_n844));
  NOR3_X1   g419(.A1(new_n832), .A2(new_n835), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT34), .B1(new_n825), .B2(new_n831), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT36), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n849), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n815), .A2(new_n851), .A3(new_n852), .ZN(G311));
  NAND3_X1  g428(.A1(new_n815), .A2(new_n851), .A3(new_n852), .ZN(G150));
  NAND2_X1  g429(.A1(new_n625), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n530), .A2(G93), .B1(G55), .B2(new_n531), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n528), .A2(G67), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n857), .B1(new_n545), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n567), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n567), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n856), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n867), .A2(new_n868), .A3(G860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n861), .A2(G860), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n869), .A2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n653), .B(KEYINPUT102), .ZN(new_n873));
  INV_X1    g448(.A(G162), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n489), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n515), .A2(new_n519), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n795), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n749), .ZN(new_n879));
  INV_X1    g454(.A(new_n765), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n503), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n468), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G142), .B2(new_n498), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n643), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n841), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(new_n880), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n881), .A2(new_n888), .A3(KEYINPUT103), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n876), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n881), .B2(new_n889), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n881), .A2(new_n888), .A3(new_n889), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n875), .B(G160), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n899), .B2(new_n892), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g478(.A1(new_n861), .A2(new_n628), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n827), .A2(G290), .ZN(new_n905));
  NAND2_X1  g480(.A1(G305), .A2(new_n614), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(G166), .A2(new_n821), .ZN(new_n908));
  NAND2_X1  g483(.A1(G303), .A2(G288), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n907), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n639), .B(new_n864), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n630), .A2(new_n624), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND2_X1  g492(.A1(G299), .A2(new_n625), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n630), .A2(KEYINPUT104), .A3(new_n624), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n916), .A2(new_n918), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n915), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n923), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n915), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n914), .B(new_n929), .Z(new_n930));
  OAI21_X1  g505(.A(new_n904), .B1(new_n930), .B2(new_n628), .ZN(G295));
  OAI21_X1  g506(.A(new_n904), .B1(new_n930), .B2(new_n628), .ZN(G331));
  AOI21_X1  g507(.A(G301), .B1(new_n591), .B2(new_n593), .ZN(new_n933));
  NOR2_X1   g508(.A1(G168), .A2(G171), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n864), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n865), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n926), .A3(new_n922), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n937), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n923), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n911), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n911), .A3(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n897), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n919), .A2(new_n921), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n938), .A2(KEYINPUT41), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n923), .B1(new_n938), .B2(new_n925), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n911), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n944), .A2(new_n951), .A3(new_n952), .A4(new_n897), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n944), .A2(new_n951), .A3(new_n897), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n957), .B2(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n944), .A2(new_n952), .A3(new_n897), .A4(new_n945), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n958), .A2(KEYINPUT107), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT107), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(G397));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n515), .B2(new_n519), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n963), .C1(new_n515), .C2(new_n519), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n480), .A2(G40), .A3(new_n488), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT46), .Z(new_n975));
  INV_X1    g550(.A(new_n749), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n795), .B(new_n797), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n979), .A2(KEYINPUT47), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(KEYINPUT47), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n749), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n841), .A2(new_n843), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n841), .A2(new_n843), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n971), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n971), .A2(new_n977), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT112), .Z(new_n990));
  NOR2_X1   g565(.A1(new_n749), .A2(new_n972), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n971), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n971), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT48), .Z(new_n996));
  OAI22_X1  g571(.A1(new_n980), .A2(new_n981), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n984), .A2(new_n986), .A3(new_n992), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n795), .A2(new_n797), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(new_n971), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1000), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT126), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n504), .A2(new_n512), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n963), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1009), .B(new_n963), .C1(new_n515), .C2(new_n519), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AND4_X1   g588(.A1(G40), .A2(new_n480), .A3(new_n753), .A4(new_n488), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n514), .B2(new_n520), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1013), .B(new_n1014), .C1(new_n1009), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  AOI211_X1 g594(.A(G1384), .B(new_n966), .C1(new_n514), .C2(new_n520), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n964), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(G40), .A3(new_n480), .A4(new_n488), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1019), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n513), .B1(new_n504), .B2(new_n512), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n515), .A2(new_n519), .A3(KEYINPUT72), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n963), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(KEYINPUT116), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1018), .A2(G168), .A3(new_n1024), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1024), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1027), .A2(KEYINPUT50), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT116), .B1(new_n1035), .B2(new_n1014), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n592), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT51), .A3(G8), .A4(new_n1030), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1033), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1006), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT119), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1033), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT62), .A3(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n970), .A2(new_n964), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n821), .A2(G1976), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1047), .A2(G8), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1048), .B(G8), .C1(new_n970), .C2(new_n964), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n602), .A2(new_n603), .ZN(new_n1055));
  INV_X1    g630(.A(new_n605), .ZN(new_n1056));
  OAI21_X1  g631(.A(G1981), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n607), .A2(new_n1058), .A3(new_n603), .A4(new_n602), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT49), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1047), .A2(G8), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1054), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT113), .B(G1971), .Z(new_n1065));
  INV_X1    g640(.A(new_n966), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n521), .B2(new_n963), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT45), .B(new_n963), .C1(new_n515), .C2(new_n519), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n480), .A3(G40), .A4(new_n488), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n970), .B1(KEYINPUT50), .B2(new_n964), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(KEYINPUT50), .B2(new_n1027), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(G2090), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n537), .A2(new_n538), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(G8), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G8), .ZN(new_n1082));
  INV_X1    g657(.A(G2090), .ZN(new_n1083));
  INV_X1    g658(.A(new_n970), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1035), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1085), .B2(new_n1070), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1079), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1086), .B2(new_n1079), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1064), .B(new_n1081), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AND4_X1   g665(.A1(G40), .A2(new_n1068), .A3(new_n480), .A4(new_n488), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n736), .C1(new_n1066), .C2(new_n1015), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT53), .A3(new_n736), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1013), .B(new_n1084), .C1(new_n1009), .C2(new_n1015), .ZN(new_n1097));
  INV_X1    g672(.A(G1961), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1042), .A2(new_n1046), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n821), .A2(new_n1049), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1059), .ZN(new_n1106));
  OAI211_X1 g681(.A(G8), .B(new_n1047), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1064), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G286), .A2(new_n1082), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1090), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1086), .A2(new_n1079), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1115), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1108), .A2(new_n1116), .A3(new_n1064), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1103), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1097), .A2(new_n787), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(G2067), .B2(new_n1047), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n625), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n582), .B2(KEYINPUT117), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G299), .B(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1072), .A2(new_n812), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT56), .B(G2072), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1124), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1134), .A2(new_n1135), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1121), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n624), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1133), .A2(KEYINPUT61), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(new_n1142), .A3(new_n1128), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1130), .A2(new_n972), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n1047), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n567), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT59), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1121), .A2(new_n1138), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1151), .A2(new_n1139), .A3(new_n624), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1137), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n736), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n468), .B1(new_n484), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n482), .A2(KEYINPUT121), .A3(new_n483), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1068), .A2(new_n480), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n969), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n969), .A2(new_n1159), .A3(KEYINPUT122), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1162), .A2(new_n1163), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1099), .A2(KEYINPUT120), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1097), .A2(new_n1166), .A3(new_n1098), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1164), .A2(new_n1165), .A3(G301), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT54), .B1(new_n1168), .B2(new_n1101), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT123), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1067), .A2(G2078), .A3(new_n1069), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n969), .A2(new_n1159), .A3(KEYINPUT122), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT122), .B1(new_n969), .B2(new_n1159), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n1171), .A2(KEYINPUT53), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1166), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(G301), .B1(new_n1176), .B2(new_n1167), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1094), .A2(new_n1096), .A3(new_n1099), .A4(G301), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT54), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT124), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1181));
  AOI21_X1  g756(.A(G1961), .B1(new_n1035), .B2(new_n1084), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1181), .B(new_n1094), .C1(new_n1182), .C2(new_n1166), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1167), .ZN(new_n1184));
  OAI21_X1  g759(.A(G171), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT54), .A4(new_n1178), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1090), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1170), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1153), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1170), .A2(new_n1188), .A3(new_n1189), .A4(KEYINPUT125), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1119), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AND2_X1   g769(.A1(G290), .A2(G1986), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n971), .B1(new_n1195), .B2(new_n994), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n984), .A2(new_n1196), .A3(new_n988), .A4(new_n992), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1005), .B1(new_n1194), .B2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g773(.A1(new_n697), .A2(new_n699), .A3(G319), .ZN(new_n1200));
  AND2_X1   g774(.A1(new_n677), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g775(.A(G229), .ZN(new_n1202));
  OAI211_X1 g776(.A(new_n1201), .B(new_n1202), .C1(new_n895), .C2(new_n900), .ZN(new_n1203));
  AOI211_X1 g777(.A(KEYINPUT127), .B(new_n1203), .C1(new_n947), .C2(new_n953), .ZN(new_n1204));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n1205));
  INV_X1    g779(.A(new_n1203), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n954), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g781(.A1(new_n1204), .A2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n954), .A2(new_n1206), .ZN(G225));
endmodule


