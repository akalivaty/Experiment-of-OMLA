

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U327 ( .A(n460), .B(n459), .ZN(n506) );
  XOR2_X1 U328 ( .A(n480), .B(KEYINPUT28), .Z(n537) );
  XOR2_X1 U329 ( .A(G190GAT), .B(G134GAT), .Z(n295) );
  XOR2_X1 U330 ( .A(n439), .B(n304), .Z(n296) );
  OR2_X1 U331 ( .A1(n523), .A2(n525), .ZN(n422) );
  OR2_X1 U332 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U333 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U334 ( .A(n435), .B(n334), .ZN(n335) );
  XNOR2_X1 U335 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n475) );
  INV_X1 U336 ( .A(G120GAT), .ZN(n308) );
  XNOR2_X1 U337 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U338 ( .A(n476), .B(n475), .ZN(n534) );
  NOR2_X1 U339 ( .A1(n587), .A2(n457), .ZN(n458) );
  XNOR2_X1 U340 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U341 ( .A(n342), .B(n341), .ZN(n346) );
  XNOR2_X1 U342 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U343 ( .A(KEYINPUT38), .B(KEYINPUT108), .ZN(n459) );
  NOR2_X1 U344 ( .A1(n525), .A2(n482), .ZN(n566) );
  INV_X1 U345 ( .A(G43GAT), .ZN(n461) );
  XNOR2_X1 U346 ( .A(n486), .B(G183GAT), .ZN(n487) );
  XNOR2_X1 U347 ( .A(n461), .B(KEYINPUT40), .ZN(n462) );
  XNOR2_X1 U348 ( .A(n488), .B(n487), .ZN(G1350GAT) );
  XNOR2_X1 U349 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT85), .B(G71GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(G176GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U353 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n300) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n313) );
  XOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .Z(n439) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(G99GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n295), .B(n303), .ZN(n304) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n296), .B(n305), .ZN(n311) );
  XOR2_X1 U362 ( .A(G183GAT), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n409) );
  XNOR2_X1 U365 ( .A(n409), .B(G127GAT), .ZN(n309) );
  XOR2_X1 U366 ( .A(n313), .B(n312), .Z(n535) );
  INV_X1 U367 ( .A(n535), .ZN(n525) );
  XOR2_X1 U368 ( .A(G43GAT), .B(G50GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n351) );
  XOR2_X1 U371 ( .A(G169GAT), .B(G8GAT), .Z(n410) );
  XOR2_X1 U372 ( .A(n351), .B(n410), .Z(n317) );
  NAND2_X1 U373 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G22GAT), .Z(n381) );
  XOR2_X1 U376 ( .A(n318), .B(n381), .Z(n320) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G36GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT68), .B(G197GAT), .Z(n322) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(G141GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U382 ( .A(KEYINPUT30), .B(G1GAT), .Z(n324) );
  XNOR2_X1 U383 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U385 ( .A(n326), .B(n325), .Z(n327) );
  XOR2_X1 U386 ( .A(n328), .B(n327), .Z(n539) );
  XOR2_X1 U387 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n330) );
  XOR2_X1 U388 ( .A(G106GAT), .B(G78GAT), .Z(n386) );
  XOR2_X1 U389 ( .A(G71GAT), .B(KEYINPUT13), .Z(n371) );
  XNOR2_X1 U390 ( .A(n386), .B(n371), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n336) );
  XNOR2_X1 U392 ( .A(G120GAT), .B(G85GAT), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n331), .B(G57GAT), .ZN(n435) );
  NAND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  INV_X1 U395 ( .A(KEYINPUT73), .ZN(n332) );
  XOR2_X1 U396 ( .A(n336), .B(n335), .Z(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n338) );
  XNOR2_X1 U398 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n340) );
  XNOR2_X1 U400 ( .A(G99GAT), .B(G148GAT), .ZN(n339) );
  XOR2_X1 U401 ( .A(G92GAT), .B(G64GAT), .Z(n344) );
  XNOR2_X1 U402 ( .A(G176GAT), .B(KEYINPUT71), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(G204GAT), .B(n345), .Z(n418) );
  XOR2_X1 U405 ( .A(n346), .B(n418), .Z(n579) );
  NOR2_X1 U406 ( .A1(n539), .A2(n579), .ZN(n493) );
  XOR2_X1 U407 ( .A(G29GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G190GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT77), .ZN(n413) );
  XNOR2_X1 U410 ( .A(n434), .B(n413), .ZN(n349) );
  AND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(n350), .B(KEYINPUT74), .Z(n353) );
  XNOR2_X1 U414 ( .A(n351), .B(KEYINPUT76), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U416 ( .A(G85GAT), .B(G218GAT), .Z(n355) );
  XNOR2_X1 U417 ( .A(G99GAT), .B(G162GAT), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U419 ( .A(n357), .B(n356), .Z(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT75), .B(KEYINPUT66), .Z(n359) );
  XNOR2_X1 U421 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U423 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n361) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U427 ( .A(n365), .B(n364), .Z(n565) );
  XOR2_X1 U428 ( .A(KEYINPUT36), .B(n565), .Z(n587) );
  XOR2_X1 U429 ( .A(G78GAT), .B(G211GAT), .Z(n367) );
  XNOR2_X1 U430 ( .A(G183GAT), .B(G155GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(G1GAT), .B(G127GAT), .Z(n432) );
  XOR2_X1 U433 ( .A(n368), .B(n432), .Z(n370) );
  XNOR2_X1 U434 ( .A(G8GAT), .B(G57GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n385) );
  XOR2_X1 U436 ( .A(KEYINPUT78), .B(n371), .Z(n373) );
  NAND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U439 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n375) );
  XNOR2_X1 U440 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U442 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U443 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n379) );
  XNOR2_X1 U444 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U448 ( .A(n385), .B(n384), .Z(n545) );
  XOR2_X1 U449 ( .A(KEYINPUT92), .B(n386), .Z(n388) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n389), .B(KEYINPUT93), .Z(n396) );
  XOR2_X1 U453 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n391) );
  XNOR2_X1 U454 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U456 ( .A(n392), .B(G155GAT), .Z(n394) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(G148GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n445) );
  XNOR2_X1 U459 ( .A(G50GAT), .B(n445), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U461 ( .A(KEYINPUT22), .B(G204GAT), .Z(n398) );
  XNOR2_X1 U462 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U464 ( .A(n400), .B(n399), .Z(n408) );
  XOR2_X1 U465 ( .A(KEYINPUT90), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U466 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U468 ( .A(G197GAT), .B(n403), .Z(n419) );
  XOR2_X1 U469 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n405) );
  XNOR2_X1 U470 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n419), .B(n406), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n480) );
  XOR2_X1 U474 ( .A(KEYINPUT100), .B(KEYINPUT78), .Z(n412) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n417) );
  XOR2_X1 U477 ( .A(n413), .B(KEYINPUT99), .Z(n415) );
  NAND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U480 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U482 ( .A(n421), .B(n420), .Z(n523) );
  XNOR2_X1 U483 ( .A(KEYINPUT103), .B(n422), .ZN(n423) );
  NOR2_X1 U484 ( .A1(n480), .A2(n423), .ZN(n425) );
  XNOR2_X1 U485 ( .A(KEYINPUT25), .B(KEYINPUT104), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U487 ( .A(n523), .B(KEYINPUT27), .Z(n451) );
  XOR2_X1 U488 ( .A(KEYINPUT26), .B(KEYINPUT102), .Z(n427) );
  NAND2_X1 U489 ( .A1(n480), .A2(n525), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n571) );
  NAND2_X1 U491 ( .A1(n451), .A2(n571), .ZN(n428) );
  NAND2_X1 U492 ( .A1(n429), .A2(n428), .ZN(n448) );
  XOR2_X1 U493 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n431) );
  XNOR2_X1 U494 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U496 ( .A(n433), .B(n432), .Z(n441) );
  XOR2_X1 U497 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n443) );
  XNOR2_X1 U503 ( .A(KEYINPUT97), .B(KEYINPUT1), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n450) );
  NAND2_X1 U507 ( .A1(n448), .A2(n450), .ZN(n449) );
  XOR2_X1 U508 ( .A(KEYINPUT105), .B(n449), .Z(n456) );
  XNOR2_X1 U509 ( .A(KEYINPUT98), .B(n450), .ZN(n521) );
  INV_X1 U510 ( .A(n451), .ZN(n452) );
  NOR2_X1 U511 ( .A1(n521), .A2(n452), .ZN(n532) );
  NAND2_X1 U512 ( .A1(n532), .A2(n537), .ZN(n453) );
  XNOR2_X1 U513 ( .A(KEYINPUT101), .B(n453), .ZN(n454) );
  NAND2_X1 U514 ( .A1(n454), .A2(n525), .ZN(n455) );
  NAND2_X1 U515 ( .A1(n456), .A2(n455), .ZN(n492) );
  NAND2_X1 U516 ( .A1(n545), .A2(n492), .ZN(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT37), .B(n458), .Z(n518) );
  NAND2_X1 U518 ( .A1(n493), .A2(n518), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n525), .A2(n506), .ZN(n463) );
  INV_X1 U520 ( .A(n579), .ZN(n470) );
  XNOR2_X1 U521 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n464) );
  XOR2_X1 U522 ( .A(n470), .B(n464), .Z(n541) );
  NOR2_X1 U523 ( .A1(n539), .A2(n541), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT46), .ZN(n467) );
  INV_X1 U525 ( .A(n565), .ZN(n550) );
  NAND2_X1 U526 ( .A1(n545), .A2(n550), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT47), .ZN(n474) );
  INV_X1 U528 ( .A(n539), .ZN(n574) );
  NOR2_X1 U529 ( .A1(n545), .A2(n587), .ZN(n469) );
  XNOR2_X1 U530 ( .A(KEYINPUT45), .B(n469), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n574), .A2(n472), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT120), .B(n523), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n534), .A2(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT54), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n521), .ZN(n573) );
  NOR2_X1 U538 ( .A1(n573), .A2(n480), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  INV_X1 U540 ( .A(n541), .ZN(n557) );
  NAND2_X1 U541 ( .A1(n566), .A2(n557), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(G176GAT), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1349GAT) );
  INV_X1 U545 ( .A(n545), .ZN(n583) );
  NAND2_X1 U546 ( .A1(n566), .A2(n583), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n486) );
  NOR2_X1 U548 ( .A1(n565), .A2(n545), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT16), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT83), .B(n490), .Z(n491) );
  AND2_X1 U551 ( .A1(n492), .A2(n491), .ZN(n509) );
  NAND2_X1 U552 ( .A1(n493), .A2(n509), .ZN(n501) );
  NOR2_X1 U553 ( .A1(n521), .A2(n501), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT34), .B(KEYINPUT106), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n496), .Z(G1324GAT) );
  NOR2_X1 U557 ( .A1(n523), .A2(n501), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1325GAT) );
  NOR2_X1 U560 ( .A1(n525), .A2(n501), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U563 ( .A1(n537), .A2(n501), .ZN(n502) );
  XOR2_X1 U564 ( .A(G22GAT), .B(n502), .Z(G1327GAT) );
  NOR2_X1 U565 ( .A1(n521), .A2(n506), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n523), .A2(n506), .ZN(n505) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n505), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n537), .A2(n506), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  NOR2_X1 U573 ( .A1(n574), .A2(n541), .ZN(n519) );
  NAND2_X1 U574 ( .A1(n519), .A2(n509), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n521), .A2(n515), .ZN(n510) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n515), .ZN(n512) );
  XOR2_X1 U579 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n515), .ZN(n513) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(n513), .Z(n514) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n537), .A2(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U587 ( .A(KEYINPUT111), .B(n520), .Z(n528) );
  NOR2_X1 U588 ( .A1(n521), .A2(n528), .ZN(n522) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n528), .ZN(n524) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n528), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(n526), .Z(n527) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U595 ( .A1(n537), .A2(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  INV_X1 U599 ( .A(n532), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n554) );
  NAND2_X1 U601 ( .A1(n554), .A2(n535), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT115), .B(n536), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n549) );
  NOR2_X1 U604 ( .A1(n539), .A2(n549), .ZN(n540) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n540), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n549), .ZN(n543) );
  XNOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n545), .A2(n549), .ZN(n547) );
  XNOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n554), .A2(n571), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT119), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n562), .A2(n574), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U623 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n583), .A2(n562), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n574), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n578) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .Z(n576) );
  INV_X1 U639 ( .A(n571), .ZN(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(n578), .B(n577), .Z(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n585), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n586) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

