//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n583, new_n584, new_n587, new_n589, new_n590, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n460), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G112), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n460), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n473), .B1(G124), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n461), .A2(new_n462), .ZN(new_n478));
  OR3_X1    g053(.A1(new_n478), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(new_n478), .B2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(KEYINPUT68), .B2(G114), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT68), .A2(G114), .ZN(new_n487));
  OAI211_X1 g062(.A(G2104), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G138), .A4(new_n460), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  XOR2_X1   g073(.A(new_n498), .B(KEYINPUT70), .Z(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n497), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G166));
  AOI22_X1  g091(.A1(new_n502), .A2(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n510), .A2(G51), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  AOI22_X1  g099(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n497), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n510), .A2(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  XOR2_X1   g105(.A(KEYINPUT72), .B(G81), .Z(new_n531));
  AOI22_X1  g106(.A1(new_n517), .A2(new_n531), .B1(new_n510), .B2(G43), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n497), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n535), .B2(KEYINPUT71), .ZN(new_n536));
  OR3_X1    g111(.A1(new_n534), .A2(KEYINPUT71), .A3(new_n497), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  INV_X1    g119(.A(G65), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n502), .B2(new_n504), .ZN(new_n546));
  AND2_X1   g121(.A1(G78), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(G651), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n517), .A2(G91), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n510), .A2(new_n550), .A3(G53), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n550), .B1(new_n510), .B2(G53), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n548), .B(new_n549), .C1(new_n551), .C2(new_n552), .ZN(G299));
  INV_X1    g128(.A(G171), .ZN(G301));
  INV_X1    g129(.A(G166), .ZN(G303));
  OAI21_X1  g130(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n505), .A2(G87), .A3(new_n512), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n510), .A2(G49), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  AOI22_X1  g134(.A1(new_n517), .A2(G86), .B1(new_n510), .B2(G48), .ZN(new_n560));
  INV_X1    g135(.A(G61), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n502), .B2(new_n504), .ZN(new_n562));
  NAND2_X1  g137(.A1(G73), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G305));
  AOI22_X1  g141(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n497), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n517), .A2(G85), .B1(new_n510), .B2(G47), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G290));
  NAND2_X1  g145(.A1(G301), .A2(G868), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n517), .A2(G92), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT10), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n505), .A2(G66), .ZN(new_n575));
  INV_X1    g150(.A(G79), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n500), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n571), .B1(new_n580), .B2(G868), .ZN(G321));
  XOR2_X1   g156(.A(G321), .B(KEYINPUT73), .Z(G284));
  INV_X1    g157(.A(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(G299), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(new_n583), .B2(G168), .ZN(G297));
  OAI21_X1  g160(.A(new_n584), .B1(new_n583), .B2(G168), .ZN(G280));
  INV_X1    g161(.A(G559), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n580), .B1(new_n587), .B2(G860), .ZN(G148));
  NAND2_X1  g163(.A1(new_n538), .A2(new_n583), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n579), .A2(G559), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(new_n583), .ZN(G323));
  XNOR2_X1  g166(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g167(.A1(new_n493), .A2(new_n467), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT12), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(G2100), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n479), .A2(new_n480), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G135), .ZN(new_n599));
  OAI21_X1  g174(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT75), .ZN(new_n601));
  INV_X1    g176(.A(G111), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n600), .A2(KEYINPUT75), .B1(new_n602), .B2(G2105), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n601), .A2(new_n603), .B1(new_n476), .B2(G123), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(G2096), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n596), .A2(G2100), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(G2096), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n597), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(G156));
  XNOR2_X1  g184(.A(KEYINPUT15), .B(G2435), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT76), .B(G2438), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(G2427), .B(G2430), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n614), .A2(KEYINPUT14), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2451), .B(G2454), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT16), .ZN(new_n618));
  XOR2_X1   g193(.A(G1341), .B(G1348), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n616), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(G2443), .B(G2446), .Z(new_n622));
  OAI21_X1  g197(.A(G14), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n621), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT77), .ZN(G401));
  INV_X1    g200(.A(KEYINPUT18), .ZN(new_n626));
  XOR2_X1   g201(.A(G2084), .B(G2090), .Z(new_n627));
  XNOR2_X1  g202(.A(G2067), .B(G2678), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT17), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n629), .B2(KEYINPUT18), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(G227));
  XOR2_X1   g212(.A(G1971), .B(G1976), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT19), .ZN(new_n639));
  XOR2_X1   g214(.A(G1956), .B(G2474), .Z(new_n640));
  XOR2_X1   g215(.A(G1961), .B(G1966), .Z(new_n641));
  AND2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT20), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n639), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n639), .B2(new_n645), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT79), .ZN(new_n651));
  XOR2_X1   g226(.A(G1981), .B(G1986), .Z(new_n652));
  XNOR2_X1  g227(.A(G1991), .B(G1996), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G229));
  XOR2_X1   g235(.A(KEYINPUT31), .B(G11), .Z(new_n661));
  INV_X1    g236(.A(G28), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(KEYINPUT30), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  AOI21_X1  g239(.A(G29), .B1(new_n662), .B2(KEYINPUT30), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G34), .ZN(new_n667));
  AOI21_X1  g242(.A(G29), .B1(new_n667), .B2(KEYINPUT24), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(KEYINPUT24), .B2(new_n667), .ZN(new_n669));
  INV_X1    g244(.A(G160), .ZN(new_n670));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G2084), .ZN(new_n673));
  OAI221_X1 g248(.A(new_n666), .B1(new_n672), .B2(new_n673), .C1(new_n605), .C2(new_n671), .ZN(new_n674));
  INV_X1    g249(.A(G2078), .ZN(new_n675));
  NOR2_X1   g250(.A1(G27), .A2(G29), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G164), .B2(G29), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G21), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G168), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT85), .B(G1966), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(G5), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G171), .B2(new_n680), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n686), .A2(G1961), .B1(G2078), .B2(new_n677), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n672), .A2(new_n673), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT87), .Z(new_n689));
  AND4_X1   g264(.A1(new_n679), .A2(new_n684), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G29), .A2(G33), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT25), .Z(new_n693));
  AOI22_X1  g268(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  INV_X1    g269(.A(G139), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n693), .B1(new_n460), .B2(new_n694), .C1(new_n481), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT84), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(G29), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G2072), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n671), .A2(G32), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n476), .A2(G129), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n467), .A2(G105), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n598), .B2(G141), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n700), .B1(new_n707), .B2(new_n671), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n700), .B(new_n709), .C1(new_n707), .C2(new_n671), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n711), .B(new_n712), .C1(G1961), .C2(new_n686), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n698), .B2(G2072), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n690), .A2(new_n699), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT88), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n690), .A2(new_n717), .A3(new_n699), .A4(new_n714), .ZN(new_n718));
  INV_X1    g293(.A(G2090), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n671), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n671), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n719), .A3(new_n723), .ZN(new_n726));
  INV_X1    g301(.A(G1341), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n680), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n538), .B2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n680), .A2(G4), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n580), .B2(new_n680), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1348), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n727), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n671), .A2(G26), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n479), .A2(G140), .A3(new_n480), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n738));
  INV_X1    g313(.A(G116), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G2105), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G128), .B2(new_n476), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n680), .A2(G20), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT23), .Z(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G299), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G1956), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR4_X1   g325(.A1(new_n730), .A2(new_n733), .A3(new_n745), .A4(new_n750), .ZN(new_n751));
  AND4_X1   g326(.A1(new_n716), .A2(new_n718), .A3(new_n725), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n680), .A2(G22), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G166), .B2(new_n680), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1971), .Z(new_n755));
  AND2_X1   g330(.A1(new_n680), .A2(G23), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G288), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT83), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT33), .B(G1976), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n755), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT81), .B(KEYINPUT34), .Z(new_n763));
  OR2_X1    g338(.A1(G6), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G305), .B2(new_n680), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(KEYINPUT82), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT32), .B(G1981), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n765), .A2(KEYINPUT82), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n769), .B1(new_n767), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n762), .A2(new_n763), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n671), .A2(G25), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n598), .A2(G131), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(G107), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G2105), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G119), .B2(new_n476), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(new_n671), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT35), .B(G1991), .Z(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n680), .A2(G24), .ZN(new_n787));
  INV_X1    g362(.A(G290), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n680), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT80), .B(G1986), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n774), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n763), .B1(new_n762), .B2(new_n773), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT36), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT36), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n796), .A2(new_n797), .A3(new_n774), .A4(new_n792), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n752), .A2(KEYINPUT90), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(KEYINPUT90), .B1(new_n752), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(G311));
  NAND2_X1  g377(.A1(new_n752), .A2(new_n799), .ZN(G150));
  XNOR2_X1  g378(.A(KEYINPUT94), .B(G860), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n587), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n497), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT92), .B(G55), .Z(new_n812));
  AOI22_X1  g387(.A1(new_n517), .A2(G93), .B1(new_n510), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n811), .B1(new_n810), .B2(new_n813), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n538), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n816), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n818), .A2(new_n537), .A3(new_n536), .A4(new_n814), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n808), .B(new_n820), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n805), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(KEYINPUT39), .B2(new_n822), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n810), .A2(new_n813), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n805), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(G145));
  INV_X1    g403(.A(new_n594), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n776), .A2(KEYINPUT97), .A3(new_n780), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT97), .B1(new_n776), .B2(new_n780), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n781), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n776), .A2(KEYINPUT97), .A3(new_n780), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n594), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n598), .A2(G142), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n476), .A2(G130), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT96), .Z(new_n839));
  OR2_X1    g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n832), .A2(new_n836), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n832), .B2(new_n836), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n707), .A2(new_n742), .ZN(new_n847));
  INV_X1    g422(.A(new_n706), .ZN(new_n848));
  INV_X1    g423(.A(G141), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n481), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n850), .A2(new_n737), .A3(new_n741), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n847), .A2(new_n851), .A3(G164), .ZN(new_n852));
  AOI21_X1  g427(.A(G164), .B1(new_n847), .B2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT84), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n696), .B(new_n854), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(KEYINPUT95), .ZN(new_n856));
  INV_X1    g431(.A(new_n853), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n847), .A2(new_n851), .A3(G164), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n696), .B1(new_n854), .B2(KEYINPUT95), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n846), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n845), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n832), .A2(new_n836), .A3(new_n843), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n867), .A2(KEYINPUT99), .A3(new_n856), .A4(new_n860), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n846), .B2(new_n861), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n846), .A2(new_n861), .A3(KEYINPUT98), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n864), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n605), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n862), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n846), .A2(new_n861), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g457(.A(G290), .B(G305), .Z(new_n883));
  XNOR2_X1  g458(.A(G166), .B(G288), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n883), .B(new_n884), .Z(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n820), .B(new_n590), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n579), .A2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n579), .A2(G299), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n891), .B(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n887), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n887), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n825), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(G868), .B2(new_n903), .ZN(G295));
  OAI21_X1  g479(.A(new_n902), .B1(G868), .B2(new_n903), .ZN(G331));
  XNOR2_X1  g480(.A(G171), .B(G168), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n817), .A2(new_n819), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n817), .B2(new_n819), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n908), .A3(new_n891), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  INV_X1    g486(.A(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n820), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT102), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n909), .B1(new_n915), .B2(new_n895), .ZN(new_n916));
  INV_X1    g491(.A(new_n885), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n907), .A2(new_n908), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n891), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(new_n891), .B2(KEYINPUT41), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n894), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n919), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n898), .A2(new_n911), .A3(new_n914), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n885), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n918), .A2(KEYINPUT43), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n896), .B1(new_n914), .B2(new_n911), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n885), .B1(new_n929), .B2(new_n909), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT43), .B1(new_n918), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n918), .A2(new_n934), .A3(new_n927), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n918), .B2(new_n930), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n937), .ZN(G397));
  XOR2_X1   g513(.A(KEYINPUT111), .B(G8), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n492), .A2(new_n495), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n488), .A2(new_n489), .ZN(new_n941));
  AOI21_X1  g516(.A(G1384), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(KEYINPUT105), .B(G40), .Z(new_n943));
  NOR3_X1   g518(.A1(new_n465), .A2(new_n469), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n939), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n517), .A2(G87), .B1(new_n510), .B2(G49), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(G1976), .A3(new_n556), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(KEYINPUT112), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(KEYINPUT52), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G1976), .B1(new_n946), .B2(new_n556), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT113), .B1(new_n953), .B2(KEYINPUT52), .ZN(new_n954));
  INV_X1    g529(.A(G1976), .ZN(new_n955));
  NAND2_X1  g530(.A1(G288), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n945), .A3(new_n959), .A4(new_n947), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n961));
  INV_X1    g536(.A(G1981), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n560), .A2(new_n962), .A3(new_n565), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n560), .B2(new_n565), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G305), .A2(G1981), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n560), .A2(new_n962), .A3(new_n565), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(KEYINPUT49), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n968), .A3(new_n945), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n952), .A2(new_n960), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(G166), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT55), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n944), .A2(new_n719), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n940), .A2(new_n941), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n975), .A2(new_n979), .A3(KEYINPUT110), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n978), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n974), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OR3_X1    g559(.A1(new_n465), .A2(new_n469), .A3(new_n943), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n976), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n988));
  AOI21_X1  g563(.A(G1971), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n973), .B(G8), .C1(new_n984), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n945), .ZN(new_n991));
  NOR2_X1   g566(.A1(G288), .A2(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n963), .B1(new_n969), .B2(new_n992), .ZN(new_n993));
  OAI22_X1  g568(.A1(new_n970), .A2(new_n990), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n986), .B1(G164), .B2(G1384), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(new_n988), .A3(new_n675), .A4(new_n944), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n675), .A2(KEYINPUT53), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n987), .A2(new_n988), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n985), .B1(new_n980), .B2(new_n983), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1000), .B(new_n1002), .C1(new_n1003), .C2(G1961), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n973), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n975), .A2(new_n979), .A3(new_n944), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  AOI21_X1  g584(.A(G2090), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n975), .A2(new_n979), .A3(KEYINPUT115), .A4(new_n944), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n989), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1007), .B1(new_n1012), .B2(new_n939), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n969), .A2(new_n960), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n958), .B1(new_n948), .B2(new_n949), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n951), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1006), .A2(new_n1013), .A3(new_n990), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G168), .A2(new_n939), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1003), .A2(new_n673), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1966), .B1(new_n987), .B2(new_n988), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n939), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g602(.A(G2084), .B(new_n985), .C1(new_n980), .C2(new_n983), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1020), .B1(new_n1029), .B2(new_n1019), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(G286), .A3(new_n1026), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1017), .B1(new_n1032), .B2(KEYINPUT62), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1027), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n971), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT51), .B1(new_n1035), .B2(new_n1018), .ZN(new_n1036));
  AOI211_X1 g611(.A(G168), .B(new_n939), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n996), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n944), .B1(new_n942), .B2(new_n977), .ZN(new_n1043));
  NOR3_X1   g618(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n749), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT56), .B(G2072), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n997), .A2(new_n988), .A3(new_n944), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1042), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n987), .A2(KEYINPUT120), .A3(new_n988), .A4(new_n1047), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1046), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(KEYINPUT121), .A4(new_n1045), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n1056));
  OAI21_X1  g631(.A(G299), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT119), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(G299), .B(new_n1059), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1051), .A2(new_n1054), .A3(new_n1064), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n1053), .A2(new_n1052), .A3(new_n1063), .A4(new_n1045), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G2067), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n942), .A2(new_n1070), .A3(new_n944), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n579), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1071), .B(new_n1073), .C1(new_n1003), .C2(G1348), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1072), .B2(new_n579), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n980), .A2(new_n983), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n944), .ZN(new_n1077));
  INV_X1    g652(.A(G1348), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(KEYINPUT60), .A3(new_n580), .A4(new_n1071), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1048), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1082), .A2(KEYINPUT120), .B1(new_n749), .B2(new_n1008), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1063), .B1(new_n1083), .B2(new_n1053), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1067), .B1(new_n1084), .B2(new_n1066), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n942), .B2(new_n944), .ZN(new_n1089));
  INV_X1    g664(.A(G1996), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n997), .A2(new_n988), .A3(new_n1090), .A4(new_n944), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n987), .A2(KEYINPUT122), .A3(new_n1090), .A4(new_n988), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1086), .B1(new_n1095), .B2(new_n539), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1098));
  AOI211_X1 g673(.A(new_n538), .B(new_n1098), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1069), .A2(new_n1081), .A3(new_n1085), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n579), .B1(new_n1079), .B2(new_n1071), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1066), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(new_n1065), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1000), .B1(new_n1003), .B2(G1961), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n988), .A2(new_n1001), .ZN(new_n1108));
  AND2_X1   g683(.A1(G160), .A2(G40), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n997), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT125), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n997), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(G171), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1961), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1077), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(G301), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1115), .A2(new_n1118), .A3(KEYINPUT54), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1114), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(G301), .A4(new_n1000), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT54), .B1(new_n1121), .B2(new_n1005), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1013), .A2(new_n990), .A3(new_n1016), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1106), .A2(new_n1124), .A3(new_n1032), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n990), .A2(KEYINPUT63), .ZN(new_n1126));
  OAI211_X1 g701(.A(G168), .B(new_n1026), .C1(new_n1028), .C2(new_n1023), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(G8), .B1(new_n984), .B2(new_n989), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1007), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1130), .A2(new_n1016), .A3(KEYINPUT116), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT116), .B1(new_n1130), .B2(new_n1016), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT117), .B(new_n1128), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1041), .A2(new_n1125), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT106), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n737), .A2(new_n1070), .A3(new_n741), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1070), .B1(new_n737), .B2(new_n741), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1144), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(KEYINPUT106), .A3(new_n1142), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n981), .A2(new_n986), .A3(new_n944), .ZN(new_n1149));
  OR3_X1    g724(.A1(new_n1148), .A2(KEYINPUT107), .A3(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n850), .B(G1996), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1149), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT107), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT108), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1150), .A2(KEYINPUT108), .A3(new_n1154), .A4(new_n1153), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n782), .A2(new_n784), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n781), .A2(new_n785), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1152), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(G290), .B(G1986), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1152), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT109), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1140), .A2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1149), .A2(G290), .A3(G1986), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  NAND4_X1  g743(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1152), .A2(new_n1090), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT46), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n850), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(new_n1149), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT127), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1171), .B(new_n1175), .C1(new_n1149), .C2(new_n1172), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT47), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1169), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1181), .A2(KEYINPUT126), .A3(new_n1142), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1182), .A2(new_n1152), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1142), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1180), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1166), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g763(.A1(new_n624), .A2(new_n458), .A3(G227), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1190), .B1(new_n657), .B2(new_n658), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n881), .B(new_n1191), .C1(new_n935), .C2(new_n936), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


