//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(KEYINPUT67), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n470), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n462), .A2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT69), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n466), .B1(new_n485), .B2(new_n487), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G124), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n490), .A2(new_n495), .ZN(G162));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n469), .B2(new_n470), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  OAI21_X1  g081(.A(G138), .B1(new_n506), .B2(KEYINPUT70), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n471), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n484), .A2(new_n510), .A3(new_n466), .A4(new_n504), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n508), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  AND2_X1   g094(.A1(G75), .A2(G543), .ZN(new_n520));
  OAI211_X1 g095(.A(KEYINPUT72), .B(G651), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G88), .B1(new_n524), .B2(G50), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n520), .B1(new_n518), .B2(G62), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n525), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AND2_X1   g106(.A1(new_n523), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n522), .A2(G543), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n533), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n532), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  OR3_X1    g116(.A1(new_n540), .A2(new_n541), .A3(new_n528), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n540), .B2(new_n528), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n523), .A2(G90), .B1(new_n524), .B2(G52), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(new_n518), .A2(new_n522), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(new_n537), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n552), .A2(new_n553), .B1(new_n528), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n518), .A2(G65), .ZN(new_n565));
  AND2_X1   g140(.A1(G78), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n523), .A2(G91), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  OAI21_X1  g145(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n518), .A2(G87), .A3(new_n522), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n522), .A2(G49), .A3(G543), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n518), .A2(G86), .A3(new_n522), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n575), .A2(new_n576), .B1(new_n524), .B2(G48), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n515), .B2(new_n517), .ZN(new_n579));
  AND2_X1   g154(.A1(G73), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(KEYINPUT77), .A3(G86), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n584), .B(G651), .C1(new_n579), .C2(new_n580), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n577), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n523), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n528), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n523), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n518), .A2(G66), .ZN(new_n594));
  INV_X1    g169(.A(G79), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n514), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(KEYINPUT78), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(KEYINPUT78), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  XNOR2_X1  g181(.A(G297), .B(KEYINPUT79), .ZN(G280));
  AOI21_X1  g182(.A(G559), .B1(new_n599), .B2(new_n600), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G860), .B2(new_n601), .ZN(G148));
  NAND2_X1  g184(.A1(new_n555), .A2(new_n604), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n608), .B2(new_n604), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g187(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g188(.A(G323), .B(new_n613), .ZN(G282));
  NAND2_X1  g189(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  NOR2_X1   g193(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n488), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n494), .A2(G123), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n620), .B1(new_n618), .B2(new_n615), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT85), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT86), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2084), .B(G2090), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n656), .B1(new_n651), .B2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(new_n655), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n657), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n675), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n676), .A2(KEYINPUT20), .A3(new_n675), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n677), .B1(new_n675), .B2(new_n673), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n668), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n667), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(new_n488), .A2(G139), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT25), .Z(new_n696));
  AOI22_X1  g271(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n696), .C1(new_n466), .C2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT97), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G33), .B(new_n702), .S(G29), .Z(new_n703));
  NOR2_X1   g278(.A1(G29), .A2(G35), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G162), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT29), .B(G2090), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n703), .A2(G2072), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G27), .A2(G29), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G164), .B2(G29), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G2078), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(G168), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G21), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n707), .B(new_n715), .C1(G2072), .C2(new_n703), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT31), .B(G11), .Z(new_n717));
  INV_X1    g292(.A(G28), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT99), .Z(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n722), .B1(new_n723), .B2(new_n625), .C1(new_n713), .C2(new_n714), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  INV_X1    g300(.A(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G160), .B2(new_n723), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G2084), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(G2084), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n724), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT91), .B(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n556), .B2(new_n733), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n723), .A2(G26), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT28), .Z(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(G116), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G2105), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n494), .B2(G128), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n488), .A2(KEYINPUT96), .A3(G140), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT96), .B1(new_n488), .B2(G140), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2067), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n711), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n711), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n732), .A2(new_n736), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT95), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n601), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1348), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n723), .A2(G32), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n494), .A2(G129), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G141), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND3_X1  g337(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(new_n723), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT101), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n733), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G299), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n711), .ZN(new_n774));
  INV_X1    g349(.A(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n768), .B(new_n776), .C1(new_n705), .C2(new_n706), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n716), .A2(new_n752), .A3(new_n756), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n733), .ZN(new_n780));
  NAND2_X1  g355(.A1(G166), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G22), .B2(new_n780), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT94), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(G1971), .A3(new_n784), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n790));
  NAND2_X1  g365(.A1(G288), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT93), .A4(new_n573), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n789), .B1(new_n793), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT33), .B(G1976), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n787), .A2(new_n788), .A3(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G6), .B(G305), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT32), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1981), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n797), .A2(new_n800), .A3(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n733), .A2(G24), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT92), .Z(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G290), .B2(new_n780), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1986), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n723), .A2(G25), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n494), .A2(G119), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n488), .A2(G131), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n466), .A2(G107), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT90), .Z(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(new_n723), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n805), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n801), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT34), .B1(new_n797), .B2(new_n800), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n779), .B1(new_n821), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n778), .ZN(G150));
  AOI22_X1  g401(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n528), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n547), .A2(new_n829), .B1(new_n537), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT102), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT102), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n835));
  OR3_X1    g410(.A1(new_n555), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  OAI211_X1 g412(.A(KEYINPUT103), .B(new_n828), .C1(new_n832), .C2(new_n833), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(new_n555), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n601), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n834), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(G164), .B(KEYINPUT104), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(new_n742), .C1(new_n744), .C2(new_n743), .ZN(new_n851));
  INV_X1    g426(.A(new_n502), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n504), .B1(new_n464), .B2(new_n510), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n471), .A2(new_n505), .A3(new_n507), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT104), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n857));
  NAND2_X1  g432(.A1(G164), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n745), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n851), .A2(new_n765), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n765), .B1(new_n851), .B2(new_n860), .ZN(new_n863));
  OAI211_X1 g438(.A(KEYINPUT105), .B(new_n702), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n494), .A2(G130), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n488), .A2(G142), .ZN(new_n866));
  OR2_X1    g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n617), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n811), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n851), .A2(new_n860), .ZN(new_n872));
  INV_X1    g447(.A(new_n765), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n700), .A2(new_n876), .A3(new_n701), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n861), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n864), .A2(new_n871), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n871), .B1(new_n864), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n625), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n879), .B2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g463(.A(new_n608), .B(new_n840), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n598), .A2(G299), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n773), .A2(new_n593), .A3(new_n597), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n893), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n793), .B(G290), .ZN(new_n900));
  XNOR2_X1  g475(.A(G305), .B(G303), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n894), .A2(new_n903), .A3(new_n897), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n899), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n899), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(G868), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n834), .A2(new_n604), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(G295));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n908), .ZN(G331));
  XNOR2_X1  g485(.A(G301), .B(G168), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n840), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n836), .A2(new_n911), .A3(new_n839), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n896), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n893), .A3(new_n914), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n902), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT106), .B1(new_n915), .B2(new_n896), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n902), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n918), .ZN(new_n925));
  INV_X1    g500(.A(new_n902), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n920), .A4(new_n919), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT44), .Z(G397));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT45), .B1(new_n850), .B2(new_n932), .ZN(new_n933));
  AND4_X1   g508(.A1(G40), .A2(new_n468), .A3(new_n475), .A4(new_n481), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(KEYINPUT107), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n934), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(G1996), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n745), .B(G2067), .Z(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n765), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n935), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(KEYINPUT125), .A3(new_n946), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT47), .A3(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n939), .A2(G1986), .A3(G290), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT48), .Z(new_n953));
  OAI21_X1  g528(.A(new_n944), .B1(new_n936), .B2(new_n765), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n941), .A2(new_n765), .B1(new_n935), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n811), .B(new_n815), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n935), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n812), .A3(new_n814), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(G2067), .B2(new_n745), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n935), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT47), .B1(new_n949), .B2(new_n950), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  AND3_X1   g540(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  NOR2_X1   g544(.A1(G164), .A2(G1384), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT110), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G2090), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n855), .A2(new_n976), .A3(new_n932), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT109), .B1(G164), .B2(G1384), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n971), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n974), .A2(new_n975), .A3(new_n934), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n856), .A2(new_n858), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n934), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n786), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n965), .B(new_n968), .C1(new_n980), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n581), .ZN(new_n989));
  INV_X1    g564(.A(G48), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n576), .B1(new_n990), .B2(new_n537), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G305), .B2(G1981), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n934), .A2(new_n977), .A3(new_n978), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n993), .A2(new_n999), .A3(new_n994), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n993), .B2(new_n994), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n995), .B(new_n998), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n793), .A2(KEYINPUT111), .A3(G1976), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n791), .A2(G1976), .A3(new_n792), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT52), .B1(new_n1007), .B2(new_n997), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n998), .A2(new_n1003), .A3(new_n1006), .A4(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G288), .A2(G1976), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1002), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n997), .B(KEYINPUT113), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n988), .A2(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1012), .A2(new_n987), .ZN(new_n1018));
  INV_X1    g593(.A(new_n986), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n976), .B1(new_n855), .B2(new_n932), .ZN(new_n1020));
  NOR3_X1   g595(.A1(G164), .A2(KEYINPUT109), .A3(G1384), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT50), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n468), .A2(new_n475), .A3(G40), .A4(new_n481), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n970), .B2(new_n971), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2090), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(KEYINPUT114), .A3(new_n1024), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n968), .B1(new_n1028), .B2(new_n965), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n977), .B2(new_n978), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n855), .A2(new_n982), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n934), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n714), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2084), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n974), .A2(new_n1036), .A3(new_n934), .A4(new_n979), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT115), .B(new_n714), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(G8), .A3(G168), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1018), .A2(new_n1029), .A3(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n980), .A2(new_n986), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n968), .B1(new_n1045), .B2(new_n965), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1018), .A2(KEYINPUT63), .A3(new_n1041), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1017), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n1049));
  XNOR2_X1  g624(.A(G299), .B(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n855), .A2(new_n971), .A3(new_n932), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n934), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n775), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n983), .A2(new_n984), .A3(new_n934), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1050), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n974), .A2(new_n934), .A3(new_n979), .ZN(new_n1059));
  INV_X1    g634(.A(G1348), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n996), .A2(G2067), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n601), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1054), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT60), .B(new_n601), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n599), .A2(new_n1069), .A3(new_n600), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1054), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1058), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n996), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1023), .A2(G1996), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n983), .A2(new_n984), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n555), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1079), .B(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1064), .A2(new_n1057), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1050), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1074), .B(new_n1082), .C1(new_n1084), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1072), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1058), .A2(KEYINPUT118), .A3(new_n1073), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n1088), .A3(new_n1087), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(KEYINPUT119), .A3(new_n1074), .A4(new_n1082), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1065), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n965), .B1(new_n1098), .B2(new_n1035), .ZN(new_n1099));
  NAND2_X1  g674(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(G168), .B2(new_n965), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1039), .B2(G8), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1097), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1039), .A2(G8), .A3(G286), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1018), .A2(new_n1029), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n985), .B2(G2078), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1112), .B(new_n1109), .C1(new_n985), .C2(G2078), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1111), .A2(new_n1113), .B1(new_n750), .B2(new_n1059), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1109), .A2(G2078), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(G301), .B(KEYINPUT54), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n983), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n476), .A2(KEYINPUT122), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n481), .A2(G40), .A3(new_n1116), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n476), .B2(KEYINPUT122), .ZN(new_n1124));
  NOR4_X1   g699(.A1(new_n933), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1125), .B2(KEYINPUT123), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1114), .B(new_n1126), .C1(KEYINPUT123), .C2(new_n1125), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1107), .A2(new_n1108), .A3(new_n1120), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1048), .B1(new_n1096), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1018), .A2(new_n1029), .A3(new_n1118), .A4(G171), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1106), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1101), .B(new_n1097), .C1(new_n1039), .C2(G8), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1102), .A2(KEYINPUT62), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1135));
  AOI211_X1 g710(.A(KEYINPUT124), .B(new_n1130), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1130), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1129), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(G290), .B(G1986), .Z(new_n1142));
  OAI211_X1 g717(.A(new_n955), .B(new_n957), .C1(new_n939), .C2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT108), .Z(new_n1144));
  OAI21_X1  g719(.A(new_n964), .B1(new_n1141), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g720(.A1(new_n663), .A2(new_n665), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n663), .A2(new_n665), .ZN(new_n1148));
  NOR3_X1   g722(.A1(new_n1147), .A2(new_n1148), .A3(new_n460), .ZN(new_n1149));
  AND3_X1   g723(.A1(new_n1149), .A2(KEYINPUT126), .A3(new_n647), .ZN(new_n1150));
  AOI21_X1  g724(.A(KEYINPUT126), .B1(new_n1149), .B2(new_n647), .ZN(new_n1151));
  OAI211_X1 g725(.A(new_n690), .B(new_n692), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n886), .B2(new_n884), .ZN(new_n1153));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  AND3_X1   g728(.A1(new_n1153), .A2(new_n930), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1153), .B2(new_n930), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1156), .ZN(G308));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n930), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n1158), .A2(KEYINPUT127), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n930), .A3(new_n1154), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1160), .ZN(G225));
endmodule


