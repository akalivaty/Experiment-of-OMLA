

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  INV_X1 U324 ( .A(n578), .ZN(n496) );
  OR2_X1 U325 ( .A1(n589), .A2(n480), .ZN(n476) );
  XNOR2_X2 U326 ( .A(n399), .B(n398), .ZN(n480) );
  XNOR2_X1 U327 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U328 ( .A(n423), .B(n395), .ZN(n396) );
  NOR2_X1 U329 ( .A1(n563), .A2(n417), .ZN(n418) );
  XNOR2_X1 U330 ( .A(n422), .B(n352), .ZN(n356) );
  XOR2_X1 U331 ( .A(n361), .B(n360), .Z(n292) );
  NOR2_X1 U332 ( .A1(n588), .A2(n510), .ZN(n406) );
  XNOR2_X1 U333 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X1 U334 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n415) );
  INV_X1 U335 ( .A(KEYINPUT83), .ZN(n350) );
  XNOR2_X1 U336 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U337 ( .A(n362), .B(n292), .ZN(n363) );
  XNOR2_X1 U338 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U339 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U340 ( .A(n305), .B(n304), .ZN(n309) );
  XNOR2_X1 U341 ( .A(n456), .B(n455), .ZN(n539) );
  XNOR2_X1 U342 ( .A(G211GAT), .B(KEYINPUT124), .ZN(n470) );
  XNOR2_X1 U343 ( .A(n473), .B(G197GAT), .ZN(n474) );
  XNOR2_X1 U344 ( .A(n471), .B(n470), .ZN(G1354GAT) );
  XNOR2_X1 U345 ( .A(n475), .B(n474), .ZN(G1352GAT) );
  XOR2_X2 U346 ( .A(G99GAT), .B(G85GAT), .Z(n388) );
  XOR2_X1 U347 ( .A(KEYINPUT9), .B(n388), .Z(n294) );
  XOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT77), .Z(n314) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(n314), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n299) );
  XOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .Z(n330) );
  INV_X1 U352 ( .A(G92GAT), .ZN(n295) );
  XOR2_X1 U353 ( .A(n330), .B(G92GAT), .Z(n297) );
  NAND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(n299), .B(n298), .Z(n305) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U358 ( .A(n424), .B(G106GAT), .ZN(n303) );
  XOR2_X1 U359 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n301) );
  XNOR2_X1 U360 ( .A(KEYINPUT75), .B(KEYINPUT10), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U362 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n307) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U365 ( .A(KEYINPUT7), .B(n308), .ZN(n384) );
  XNOR2_X1 U366 ( .A(n309), .B(n384), .ZN(n578) );
  XOR2_X1 U367 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n311) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n319) );
  XOR2_X1 U370 ( .A(G85GAT), .B(G148GAT), .Z(n313) );
  XNOR2_X1 U371 ( .A(G127GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n315) );
  XOR2_X1 U373 ( .A(n315), .B(n314), .Z(n317) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(G162GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT4), .B(G57GAT), .Z(n321) );
  NAND2_X1 U378 ( .A1(G225GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(n322), .B(KEYINPUT95), .Z(n327) );
  XOR2_X1 U381 ( .A(G120GAT), .B(KEYINPUT85), .Z(n324) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n442) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n325), .B(KEYINPUT2), .ZN(n428) );
  XNOR2_X1 U386 ( .A(n442), .B(n428), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n563) );
  XOR2_X1 U389 ( .A(KEYINPUT96), .B(n330), .Z(n332) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n338) );
  NAND2_X1 U392 ( .A1(n295), .A2(G64GAT), .ZN(n335) );
  INV_X1 U393 ( .A(G64GAT), .ZN(n333) );
  NAND2_X1 U394 ( .A1(n333), .A2(G92GAT), .ZN(n334) );
  NAND2_X1 U395 ( .A1(n335), .A2(n334), .ZN(n337) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n389) );
  XOR2_X1 U398 ( .A(n338), .B(n389), .Z(n344) );
  XOR2_X1 U399 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n421) );
  XOR2_X1 U402 ( .A(KEYINPUT78), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n359) );
  XNOR2_X1 U405 ( .A(n421), .B(n359), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U407 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n346) );
  XNOR2_X1 U408 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(n347), .ZN(n441) );
  XOR2_X1 U411 ( .A(n348), .B(n441), .Z(n537) );
  INV_X1 U412 ( .A(n537), .ZN(n484) );
  XNOR2_X1 U413 ( .A(n484), .B(KEYINPUT119), .ZN(n414) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G155GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n349), .B(G78GAT), .ZN(n422) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XOR2_X1 U417 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n354) );
  XNOR2_X1 U418 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n358) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(G57GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n392) );
  XNOR2_X1 U424 ( .A(n359), .B(n392), .ZN(n362) );
  XOR2_X1 U425 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n361) );
  XNOR2_X1 U426 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n360) );
  XOR2_X1 U427 ( .A(G1GAT), .B(KEYINPUT70), .Z(n378) );
  XOR2_X1 U428 ( .A(G15GAT), .B(G127GAT), .Z(n450) );
  XNOR2_X1 U429 ( .A(n378), .B(n450), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n574) );
  XOR2_X1 U431 ( .A(KEYINPUT107), .B(n574), .Z(n583) );
  XOR2_X1 U432 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n368) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n382) );
  XOR2_X1 U435 ( .A(G22GAT), .B(G141GAT), .Z(n370) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(G50GAT), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U438 ( .A(G113GAT), .B(G15GAT), .Z(n372) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(G197GAT), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U441 ( .A(n374), .B(n373), .Z(n380) );
  XOR2_X1 U442 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n376) );
  NAND2_X1 U443 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U447 ( .A(n382), .B(n381), .Z(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n580) );
  INV_X1 U449 ( .A(n580), .ZN(n566) );
  XNOR2_X1 U450 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n400) );
  XOR2_X1 U451 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n386) );
  XNOR2_X1 U452 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n385) );
  XOR2_X1 U453 ( .A(n386), .B(n385), .Z(n399) );
  AND2_X1 U454 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U456 ( .A(KEYINPUT72), .B(n391), .Z(n394) );
  XNOR2_X1 U457 ( .A(n392), .B(KEYINPUT73), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n397) );
  XOR2_X1 U459 ( .A(G106GAT), .B(G148GAT), .Z(n423) );
  XOR2_X1 U460 ( .A(G120GAT), .B(G78GAT), .Z(n395) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n400), .B(n480), .ZN(n460) );
  AND2_X1 U463 ( .A1(n566), .A2(n460), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n401), .B(KEYINPUT46), .ZN(n402) );
  NOR2_X1 U465 ( .A1(n583), .A2(n402), .ZN(n403) );
  XNOR2_X1 U466 ( .A(KEYINPUT108), .B(n403), .ZN(n404) );
  AND2_X1 U467 ( .A1(n404), .A2(n496), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n405), .B(KEYINPUT47), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n496), .B(KEYINPUT36), .ZN(n588) );
  INV_X1 U470 ( .A(n574), .ZN(n510) );
  XNOR2_X1 U471 ( .A(n406), .B(KEYINPUT45), .ZN(n407) );
  NAND2_X1 U472 ( .A1(n407), .A2(n480), .ZN(n408) );
  NOR2_X1 U473 ( .A1(n566), .A2(n408), .ZN(n409) );
  XNOR2_X1 U474 ( .A(KEYINPUT109), .B(n409), .ZN(n410) );
  NAND2_X1 U475 ( .A1(n411), .A2(n410), .ZN(n413) );
  XNOR2_X1 U476 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n412) );
  XNOR2_X2 U477 ( .A(n413), .B(n412), .ZN(n546) );
  NAND2_X1 U478 ( .A1(n414), .A2(n546), .ZN(n416) );
  XOR2_X1 U479 ( .A(KEYINPUT65), .B(n418), .Z(n468) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n420) );
  XNOR2_X1 U481 ( .A(G211GAT), .B(KEYINPUT22), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n437) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n435) );
  XOR2_X1 U484 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n426) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(n427), .B(KEYINPUT93), .Z(n433) );
  INV_X1 U488 ( .A(G204GAT), .ZN(n479) );
  XOR2_X1 U489 ( .A(G204GAT), .B(n428), .Z(n430) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n431), .B(KEYINPUT90), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n486) );
  NAND2_X1 U496 ( .A1(n468), .A2(n486), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n438), .B(KEYINPUT55), .ZN(n457) );
  XOR2_X1 U498 ( .A(G183GAT), .B(KEYINPUT86), .Z(n440) );
  XNOR2_X1 U499 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n456) );
  INV_X1 U501 ( .A(n441), .ZN(n446) );
  XOR2_X1 U502 ( .A(G176GAT), .B(n442), .Z(n444) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT89), .B(G71GAT), .Z(n448) );
  XNOR2_X1 U507 ( .A(G190GAT), .B(G134GAT), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U509 ( .A(n449), .B(G99GAT), .Z(n452) );
  XNOR2_X1 U510 ( .A(G43GAT), .B(n450), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n457), .A2(n539), .ZN(n461) );
  INV_X1 U514 ( .A(n461), .ZN(n584) );
  NAND2_X1 U515 ( .A1(n578), .A2(n584), .ZN(n459) );
  XNOR2_X1 U516 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  BUF_X1 U518 ( .A(n460), .Z(n570) );
  INV_X1 U519 ( .A(n570), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n462), .A2(n461), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(G176GAT), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  NOR2_X1 U524 ( .A1(n539), .A2(n486), .ZN(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n490) );
  NAND2_X1 U527 ( .A1(n490), .A2(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT122), .B(n469), .ZN(n589) );
  INV_X1 U529 ( .A(n589), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n472), .A2(n574), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n472), .A2(n566), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n479), .B(n478), .ZN(G1353GAT) );
  NAND2_X1 U536 ( .A1(n480), .A2(n566), .ZN(n513) );
  XOR2_X1 U537 ( .A(n484), .B(KEYINPUT27), .Z(n489) );
  INV_X1 U538 ( .A(n489), .ZN(n482) );
  XNOR2_X1 U539 ( .A(KEYINPUT28), .B(n486), .ZN(n506) );
  NAND2_X1 U540 ( .A1(n563), .A2(n506), .ZN(n481) );
  NOR2_X1 U541 ( .A1(n482), .A2(n481), .ZN(n547) );
  XNOR2_X1 U542 ( .A(KEYINPUT97), .B(n547), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n539), .A2(n483), .ZN(n495) );
  INV_X1 U544 ( .A(n539), .ZN(n549) );
  NOR2_X1 U545 ( .A1(n549), .A2(n484), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(n485), .Z(n487) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT25), .B(n488), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n565) );
  XNOR2_X1 U550 ( .A(KEYINPUT99), .B(n565), .ZN(n491) );
  NOR2_X1 U551 ( .A1(n492), .A2(n491), .ZN(n493) );
  NOR2_X1 U552 ( .A1(n563), .A2(n493), .ZN(n494) );
  NOR2_X1 U553 ( .A1(n495), .A2(n494), .ZN(n509) );
  NAND2_X1 U554 ( .A1(n574), .A2(n496), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT84), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(KEYINPUT16), .ZN(n499) );
  OR2_X1 U557 ( .A1(n509), .A2(n499), .ZN(n524) );
  NOR2_X1 U558 ( .A1(n513), .A2(n524), .ZN(n507) );
  NAND2_X1 U559 ( .A1(n563), .A2(n507), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT34), .B(n500), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U562 ( .A1(n537), .A2(n507), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n504) );
  NAND2_X1 U565 ( .A1(n507), .A2(n539), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U567 ( .A(G15GAT), .B(n505), .Z(G1326GAT) );
  INV_X1 U568 ( .A(n506), .ZN(n541) );
  NAND2_X1 U569 ( .A1(n541), .A2(n507), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U571 ( .A1(n509), .A2(n588), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U573 ( .A(KEYINPUT37), .B(n512), .Z(n535) );
  NOR2_X1 U574 ( .A1(n535), .A2(n513), .ZN(n514) );
  XNOR2_X1 U575 ( .A(KEYINPUT38), .B(n514), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n563), .A2(n520), .ZN(n516) );
  XOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT39), .Z(n515) );
  XNOR2_X1 U578 ( .A(n516), .B(n515), .ZN(G1328GAT) );
  NAND2_X1 U579 ( .A1(n520), .A2(n537), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n517), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U581 ( .A1(n520), .A2(n539), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT40), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G43GAT), .B(n519), .ZN(G1330GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n541), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n523) );
  XNOR2_X1 U587 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n580), .A2(n570), .ZN(n534) );
  OR2_X1 U590 ( .A1(n524), .A2(n534), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT103), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n530), .A2(n563), .ZN(n526) );
  XOR2_X1 U593 ( .A(n527), .B(n526), .Z(G1332GAT) );
  NAND2_X1 U594 ( .A1(n537), .A2(n530), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n528), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U596 ( .A1(n539), .A2(n530), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n529), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n532) );
  NAND2_X1 U599 ( .A1(n530), .A2(n541), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U601 ( .A(G78GAT), .B(n533), .Z(G1335GAT) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n563), .A2(n542), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G85GAT), .B(n536), .ZN(G1336GAT) );
  NAND2_X1 U605 ( .A1(n537), .A2(n542), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n538), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U607 ( .A1(n539), .A2(n542), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n540), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(G106GAT), .B(n545), .Z(G1339GAT) );
  XOR2_X1 U613 ( .A(G113GAT), .B(KEYINPUT111), .Z(n551) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n560), .A2(n566), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1340GAT) );
  XOR2_X1 U618 ( .A(G120GAT), .B(KEYINPUT112), .Z(n553) );
  NAND2_X1 U619 ( .A1(n560), .A2(n570), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1341GAT) );
  XNOR2_X1 U623 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n557) );
  NAND2_X1 U625 ( .A1(n560), .A2(n583), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1342GAT) );
  XOR2_X1 U628 ( .A(G134GAT), .B(KEYINPUT51), .Z(n562) );
  NAND2_X1 U629 ( .A1(n560), .A2(n578), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1343GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n568) );
  NAND2_X1 U632 ( .A1(n563), .A2(n546), .ZN(n564) );
  NOR2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G141GAT), .B(n569), .ZN(G1344GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n572) );
  NAND2_X1 U638 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G148GAT), .B(n573), .ZN(G1345GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT118), .ZN(n576) );
  XNOR2_X1 U643 ( .A(G155GAT), .B(n576), .ZN(G1346GAT) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U646 ( .A1(n461), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1348GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n587) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U655 ( .A(n591), .B(n590), .Z(G1355GAT) );
endmodule

