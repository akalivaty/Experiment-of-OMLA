

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U321 ( .A1(n459), .A2(n446), .ZN(n564) );
  XOR2_X1 U322 ( .A(n289), .B(n344), .Z(n521) );
  XOR2_X1 U323 ( .A(KEYINPUT90), .B(n471), .Z(n519) );
  XNOR2_X1 U324 ( .A(n342), .B(n341), .ZN(n289) );
  XOR2_X1 U325 ( .A(G92GAT), .B(G218GAT), .Z(n290) );
  XNOR2_X1 U326 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n457) );
  INV_X1 U327 ( .A(KEYINPUT91), .ZN(n333) );
  XNOR2_X1 U328 ( .A(n421), .B(KEYINPUT119), .ZN(n422) );
  XNOR2_X1 U329 ( .A(n521), .B(n457), .ZN(n467) );
  XNOR2_X1 U330 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U331 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U332 ( .A(n345), .B(n335), .ZN(n337) );
  XNOR2_X1 U333 ( .A(n353), .B(n352), .ZN(n354) );
  OR2_X1 U334 ( .A1(n460), .A2(n532), .ZN(n473) );
  XNOR2_X1 U335 ( .A(n355), .B(n354), .ZN(n356) );
  INV_X1 U336 ( .A(KEYINPUT37), .ZN(n490) );
  XOR2_X1 U337 ( .A(n310), .B(n309), .Z(n532) );
  XOR2_X1 U338 ( .A(n464), .B(KEYINPUT28), .Z(n534) );
  XNOR2_X1 U339 ( .A(n451), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U340 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT65), .B(KEYINPUT20), .Z(n292) );
  XNOR2_X1 U342 ( .A(G120GAT), .B(KEYINPUT80), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U344 ( .A(G190GAT), .B(G127GAT), .Z(n294) );
  XOR2_X1 U345 ( .A(G113GAT), .B(KEYINPUT0), .Z(n316) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(n316), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U348 ( .A(n296), .B(n295), .Z(n298) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U351 ( .A(G71GAT), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U354 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT79), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(n305), .ZN(n343) );
  XOR2_X1 U359 ( .A(G176GAT), .B(G183GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(n343), .B(n308), .Z(n309) );
  INV_X1 U363 ( .A(n532), .ZN(n459) );
  XOR2_X1 U364 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n445) );
  XNOR2_X1 U365 ( .A(G1GAT), .B(G127GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n311), .B(G155GAT), .ZN(n358) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G57GAT), .Z(n385) );
  XOR2_X1 U368 ( .A(n358), .B(n385), .Z(n318) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n312), .B(G85GAT), .ZN(n349) );
  XOR2_X1 U371 ( .A(KEYINPUT1), .B(n349), .Z(n314) );
  NAND2_X1 U372 ( .A1(G225GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n320) );
  XNOR2_X1 U377 ( .A(G162GAT), .B(KEYINPUT5), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U379 ( .A(n322), .B(n321), .Z(n331) );
  XOR2_X1 U380 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n324) );
  XNOR2_X1 U381 ( .A(KEYINPUT3), .B(G148GAT), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(G141GAT), .B(n325), .Z(n442) );
  INV_X1 U384 ( .A(n442), .ZN(n329) );
  XOR2_X1 U385 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n327) );
  XNOR2_X1 U386 ( .A(KEYINPUT6), .B(KEYINPUT86), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U388 ( .A(n329), .B(n328), .Z(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n471) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n290), .B(n332), .ZN(n345) );
  NAND2_X1 U392 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n336), .B(KEYINPUT74), .ZN(n362) );
  XOR2_X1 U395 ( .A(n337), .B(n362), .Z(n342) );
  XOR2_X1 U396 ( .A(G211GAT), .B(KEYINPUT21), .Z(n339) );
  XNOR2_X1 U397 ( .A(G197GAT), .B(KEYINPUT83), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n438) );
  XNOR2_X1 U399 ( .A(G176GAT), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n340), .B(G64GAT), .ZN(n377) );
  XNOR2_X1 U401 ( .A(n438), .B(n377), .ZN(n341) );
  INV_X1 U402 ( .A(n343), .ZN(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT118), .B(n521), .ZN(n420) );
  INV_X1 U404 ( .A(KEYINPUT45), .ZN(n374) );
  XOR2_X1 U405 ( .A(G50GAT), .B(G162GAT), .Z(n439) );
  XOR2_X1 U406 ( .A(G99GAT), .B(G106GAT), .Z(n386) );
  XNOR2_X1 U407 ( .A(n439), .B(n386), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n345), .B(KEYINPUT11), .ZN(n347) );
  AND2_X1 U409 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n355) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n348), .B(KEYINPUT7), .ZN(n396) );
  XNOR2_X1 U413 ( .A(n396), .B(n349), .ZN(n353) );
  XOR2_X1 U414 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n351) );
  XNOR2_X1 U415 ( .A(KEYINPUT72), .B(KEYINPUT10), .ZN(n350) );
  XOR2_X1 U416 ( .A(n351), .B(n350), .Z(n352) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n559) );
  XOR2_X1 U418 ( .A(KEYINPUT73), .B(n559), .Z(n474) );
  INV_X1 U419 ( .A(n474), .ZN(n541) );
  XOR2_X1 U420 ( .A(n541), .B(KEYINPUT36), .Z(n581) );
  XOR2_X1 U421 ( .A(n358), .B(KEYINPUT75), .Z(n360) );
  NAND2_X1 U422 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U424 ( .A(n362), .B(n361), .Z(n364) );
  XOR2_X1 U425 ( .A(G22GAT), .B(G15GAT), .Z(n395) );
  XOR2_X1 U426 ( .A(G71GAT), .B(KEYINPUT13), .Z(n381) );
  XNOR2_X1 U427 ( .A(n395), .B(n381), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n372) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G57GAT), .Z(n366) );
  XNOR2_X1 U430 ( .A(G211GAT), .B(G78GAT), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U432 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n368) );
  XNOR2_X1 U433 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U435 ( .A(n370), .B(n369), .Z(n371) );
  XOR2_X1 U436 ( .A(n372), .B(n371), .Z(n577) );
  INV_X1 U437 ( .A(n577), .ZN(n555) );
  NOR2_X1 U438 ( .A1(n581), .A2(n555), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n392) );
  XOR2_X1 U440 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n376) );
  XNOR2_X1 U441 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U444 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U447 ( .A(G85GAT), .B(G92GAT), .Z(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n391) );
  XOR2_X1 U449 ( .A(KEYINPUT69), .B(G78GAT), .Z(n436) );
  XOR2_X1 U450 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n436), .B(n389), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n573) );
  NOR2_X1 U455 ( .A1(n392), .A2(n573), .ZN(n410) );
  XOR2_X1 U456 ( .A(G113GAT), .B(G141GAT), .Z(n394) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(G197GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n409) );
  XOR2_X1 U459 ( .A(n395), .B(G50GAT), .Z(n398) );
  XNOR2_X1 U460 ( .A(G36GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U462 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n400) );
  NAND2_X1 U463 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(n402), .B(n401), .Z(n407) );
  XOR2_X1 U466 ( .A(KEYINPUT29), .B(G8GAT), .Z(n404) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(G1GAT), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n405), .B(KEYINPUT30), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n569) );
  INV_X1 U472 ( .A(n569), .ZN(n546) );
  NAND2_X1 U473 ( .A1(n410), .A2(n546), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n416) );
  XNOR2_X1 U475 ( .A(n573), .B(KEYINPUT64), .ZN(n411) );
  XOR2_X1 U476 ( .A(n411), .B(KEYINPUT41), .Z(n536) );
  AND2_X1 U477 ( .A1(n536), .A2(n569), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n412), .B(KEYINPUT46), .ZN(n413) );
  XOR2_X1 U479 ( .A(KEYINPUT109), .B(n577), .Z(n563) );
  NOR2_X1 U480 ( .A1(n413), .A2(n563), .ZN(n414) );
  NAND2_X1 U481 ( .A1(n414), .A2(n559), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n416), .B(n415), .ZN(n417) );
  NAND2_X1 U483 ( .A1(n418), .A2(n417), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n419), .B(KEYINPUT48), .ZN(n530) );
  NAND2_X1 U485 ( .A1(n420), .A2(n530), .ZN(n423) );
  INV_X1 U486 ( .A(KEYINPUT54), .ZN(n421) );
  NOR2_X1 U487 ( .A1(n519), .A2(n424), .ZN(n567) );
  XOR2_X1 U488 ( .A(G155GAT), .B(KEYINPUT23), .Z(n426) );
  XNOR2_X1 U489 ( .A(G218GAT), .B(G106GAT), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U491 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n428) );
  XNOR2_X1 U492 ( .A(G22GAT), .B(KEYINPUT82), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U494 ( .A(n430), .B(n429), .Z(n435) );
  XOR2_X1 U495 ( .A(KEYINPUT85), .B(G204GAT), .Z(n432) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U498 ( .A(KEYINPUT24), .B(n433), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U500 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U503 ( .A(n443), .B(n442), .Z(n464) );
  NAND2_X1 U504 ( .A1(n567), .A2(n464), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U506 ( .A1(n564), .A2(n536), .ZN(n450) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .Z(n448) );
  XNOR2_X1 U508 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  NAND2_X1 U511 ( .A1(n564), .A2(n541), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n451) );
  INV_X1 U513 ( .A(G169GAT), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n569), .A2(n564), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n454), .B(KEYINPUT121), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(G1348GAT) );
  NOR2_X1 U517 ( .A1(n546), .A2(n573), .ZN(n492) );
  NAND2_X1 U518 ( .A1(n519), .A2(n467), .ZN(n528) );
  NOR2_X1 U519 ( .A1(n534), .A2(n528), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n458), .B(KEYINPUT93), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n532), .A2(n521), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n461), .A2(n464), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT95), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n464), .A2(n532), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n466), .B(n465), .ZN(n566) );
  NAND2_X1 U528 ( .A1(n467), .A2(n566), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n487) );
  NAND2_X1 U532 ( .A1(n577), .A2(n474), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  AND2_X1 U534 ( .A1(n487), .A2(n476), .ZN(n505) );
  AND2_X1 U535 ( .A1(n492), .A2(n505), .ZN(n485) );
  NAND2_X1 U536 ( .A1(n485), .A2(n519), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n478) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n485), .A2(n521), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U544 ( .A1(n485), .A2(n532), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n485), .A2(n534), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n555), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(n488), .ZN(n489) );
  NOR2_X1 U551 ( .A1(n581), .A2(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n518) );
  NAND2_X1 U553 ( .A1(n518), .A2(n492), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n493), .Z(n503) );
  NAND2_X1 U555 ( .A1(n503), .A2(n519), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT101), .Z(n498) );
  NAND2_X1 U560 ( .A1(n521), .A2(n503), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n502) );
  NAND2_X1 U563 ( .A1(n503), .A2(n532), .ZN(n500) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U567 ( .A1(n503), .A2(n534), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n508) );
  INV_X1 U570 ( .A(n536), .ZN(n549) );
  NOR2_X1 U571 ( .A1(n549), .A2(n569), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n517), .A2(n505), .ZN(n506) );
  XOR2_X1 U573 ( .A(KEYINPUT104), .B(n506), .Z(n513) );
  NAND2_X1 U574 ( .A1(n519), .A2(n513), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n521), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(KEYINPUT106), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n532), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U583 ( .A1(n534), .A2(n513), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U585 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  AND2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n525) );
  NAND2_X1 U587 ( .A1(n519), .A2(n525), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n521), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n532), .A2(n525), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n523), .B(KEYINPUT108), .ZN(n524) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U594 ( .A1(n525), .A2(n534), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  INV_X1 U597 ( .A(n528), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT111), .B(n531), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n545), .A2(n532), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n542), .A2(n569), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U605 ( .A1(n542), .A2(n536), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n542), .A2(n563), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n566), .A2(n545), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n546), .A2(n558), .ZN(n547) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n547), .Z(n548) );
  XNOR2_X1 U616 ( .A(KEYINPUT112), .B(n548), .ZN(G1344GAT) );
  NOR2_X1 U617 ( .A1(n549), .A2(n558), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT114), .B(KEYINPUT53), .Z(n551) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U621 ( .A(KEYINPUT113), .B(n552), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n558), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT115), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT124), .B(n568), .ZN(n580) );
  INV_X1 U635 ( .A(n580), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n576), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G218GAT), .B(n584), .Z(G1355GAT) );
endmodule

