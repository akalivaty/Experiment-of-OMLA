

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U557 ( .A(n754), .ZN(n752) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n535), .ZN(n907) );
  INV_X2 U559 ( .A(n707), .ZN(n754) );
  XNOR2_X2 U560 ( .A(KEYINPUT64), .B(n699), .ZN(n707) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  OR2_X1 U562 ( .A1(n722), .A2(n990), .ZN(n522) );
  OR2_X1 U563 ( .A1(n799), .A2(n798), .ZN(n523) );
  INV_X1 U564 ( .A(KEYINPUT27), .ZN(n701) );
  XNOR2_X1 U565 ( .A(n701), .B(KEYINPUT93), .ZN(n702) );
  XNOR2_X1 U566 ( .A(n703), .B(n702), .ZN(n705) );
  INV_X1 U567 ( .A(KEYINPUT30), .ZN(n735) );
  XNOR2_X1 U568 ( .A(n735), .B(KEYINPUT95), .ZN(n736) );
  NOR2_X1 U569 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U570 ( .A1(n754), .A2(G2084), .ZN(n733) );
  NOR2_X1 U571 ( .A1(G164), .A2(G1384), .ZN(n698) );
  NAND2_X1 U572 ( .A1(n902), .A2(G138), .ZN(n530) );
  INV_X1 U573 ( .A(n842), .ZN(n832) );
  INV_X1 U574 ( .A(KEYINPUT88), .ZN(n531) );
  INV_X1 U575 ( .A(KEYINPUT17), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n833), .A2(n832), .ZN(n834) );
  INV_X1 U577 ( .A(G2104), .ZN(n527) );
  INV_X1 U578 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U579 ( .A1(n527), .A2(n535), .ZN(n906) );
  NAND2_X1 U580 ( .A1(n906), .A2(G114), .ZN(n524) );
  XNOR2_X1 U581 ( .A(n524), .B(KEYINPUT86), .ZN(n534) );
  XNOR2_X2 U582 ( .A(n526), .B(n525), .ZN(n902) );
  NOR2_X4 U583 ( .A1(n527), .A2(G2105), .ZN(n903) );
  NAND2_X1 U584 ( .A1(n903), .A2(G102), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT87), .B(n528), .Z(n529) );
  NAND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U587 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U589 ( .A1(G126), .A2(n907), .ZN(n536) );
  XNOR2_X1 U590 ( .A(KEYINPUT85), .B(n536), .ZN(n537) );
  NOR2_X2 U591 ( .A1(n538), .A2(n537), .ZN(G164) );
  XOR2_X1 U592 ( .A(G2438), .B(G2454), .Z(n540) );
  XNOR2_X1 U593 ( .A(G2435), .B(G2430), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U595 ( .A(n541), .B(KEYINPUT104), .Z(n543) );
  XNOR2_X1 U596 ( .A(G1341), .B(G1348), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U598 ( .A(G2427), .B(G2443), .Z(n545) );
  XNOR2_X1 U599 ( .A(G2451), .B(G2446), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(n547), .B(n546), .Z(n548) );
  AND2_X1 U602 ( .A1(G14), .A2(n548), .ZN(G401) );
  INV_X1 U603 ( .A(G651), .ZN(n553) );
  NOR2_X1 U604 ( .A1(G543), .A2(n553), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n549), .Z(n668) );
  NAND2_X1 U606 ( .A1(G64), .A2(n668), .ZN(n552) );
  XOR2_X1 U607 ( .A(G543), .B(KEYINPUT0), .Z(n669) );
  NOR2_X1 U608 ( .A1(G651), .A2(n669), .ZN(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT68), .B(n550), .ZN(n663) );
  NAND2_X1 U610 ( .A1(G52), .A2(n663), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n560) );
  NOR2_X1 U612 ( .A1(n669), .A2(n553), .ZN(n657) );
  NAND2_X1 U613 ( .A1(n657), .A2(G77), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n554), .B(KEYINPUT72), .ZN(n557) );
  NOR2_X1 U615 ( .A1(G651), .A2(G543), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT67), .B(n555), .Z(n654) );
  NAND2_X1 U617 ( .A1(G90), .A2(n654), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U620 ( .A1(n560), .A2(n559), .ZN(G171) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U622 ( .A1(G111), .A2(n906), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G135), .A2(n902), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G123), .A2(n907), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT81), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n564), .B(KEYINPUT18), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n903), .A2(G99), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n941) );
  XNOR2_X1 U631 ( .A(G2096), .B(n941), .ZN(n569) );
  OR2_X1 U632 ( .A1(G2100), .A2(n569), .ZN(G156) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G82), .ZN(G220) );
  NAND2_X1 U636 ( .A1(G88), .A2(n654), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G75), .A2(n657), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G50), .A2(n663), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n668), .A2(G62), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U642 ( .A1(n575), .A2(n574), .ZN(G166) );
  NAND2_X1 U643 ( .A1(G101), .A2(n903), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(KEYINPUT69), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT23), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G113), .A2(n906), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G125), .A2(n907), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G137), .A2(n902), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n583), .A2(n582), .ZN(G160) );
  XOR2_X1 U652 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n585) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n585), .B(n584), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n851) );
  NAND2_X1 U656 ( .A1(n851), .A2(G567), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  NAND2_X1 U658 ( .A1(n668), .A2(G56), .ZN(n587) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n587), .Z(n593) );
  NAND2_X1 U660 ( .A1(n654), .A2(G81), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G68), .A2(n657), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(n591), .Z(n592) );
  NOR2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT74), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G43), .A2(n663), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n1004) );
  INV_X1 U669 ( .A(G860), .ZN(n638) );
  OR2_X1 U670 ( .A1(n1004), .A2(n638), .ZN(G153) );
  INV_X1 U671 ( .A(G868), .ZN(n627) );
  NOR2_X1 U672 ( .A1(n627), .A2(G171), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT75), .ZN(n608) );
  NAND2_X1 U674 ( .A1(G66), .A2(n668), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT76), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G92), .A2(n654), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G54), .A2(n663), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G79), .A2(n657), .ZN(n601) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(n601), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n606), .Z(n990) );
  NAND2_X1 U684 ( .A1(n627), .A2(n990), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G284) );
  NAND2_X1 U686 ( .A1(G51), .A2(n663), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT78), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G63), .A2(n668), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U690 ( .A(KEYINPUT6), .B(n612), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n654), .A2(G89), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT4), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G76), .A2(n657), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U695 ( .A(n616), .B(KEYINPUT5), .Z(n617) );
  NOR2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT79), .B(n619), .Z(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT7), .B(n620), .Z(G168) );
  XOR2_X1 U699 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U700 ( .A1(G65), .A2(n668), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G53), .A2(n663), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G91), .A2(n654), .ZN(n624) );
  NAND2_X1 U704 ( .A1(G78), .A2(n657), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n987) );
  INV_X1 U707 ( .A(n987), .ZN(G299) );
  NOR2_X1 U708 ( .A1(G286), .A2(n627), .ZN(n629) );
  NOR2_X1 U709 ( .A1(G868), .A2(G299), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U711 ( .A(KEYINPUT80), .B(n630), .ZN(G297) );
  NAND2_X1 U712 ( .A1(n638), .A2(G559), .ZN(n631) );
  INV_X1 U713 ( .A(n990), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n631), .A2(n636), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U716 ( .A1(G868), .A2(n1004), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G868), .A2(n636), .ZN(n633) );
  NOR2_X1 U718 ( .A1(G559), .A2(n633), .ZN(n634) );
  NOR2_X1 U719 ( .A1(n635), .A2(n634), .ZN(G282) );
  NAND2_X1 U720 ( .A1(G559), .A2(n636), .ZN(n637) );
  XOR2_X1 U721 ( .A(n1004), .B(n637), .Z(n677) );
  NAND2_X1 U722 ( .A1(n638), .A2(n677), .ZN(n645) );
  NAND2_X1 U723 ( .A1(G67), .A2(n668), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G55), .A2(n663), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G93), .A2(n654), .ZN(n642) );
  NAND2_X1 U727 ( .A1(G80), .A2(n657), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n679) );
  XOR2_X1 U730 ( .A(n645), .B(n679), .Z(G145) );
  NAND2_X1 U731 ( .A1(G85), .A2(n654), .ZN(n646) );
  XNOR2_X1 U732 ( .A(n646), .B(KEYINPUT70), .ZN(n653) );
  NAND2_X1 U733 ( .A1(G72), .A2(n657), .ZN(n648) );
  NAND2_X1 U734 ( .A1(G60), .A2(n668), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U736 ( .A1(G47), .A2(n663), .ZN(n649) );
  XNOR2_X1 U737 ( .A(KEYINPUT71), .B(n649), .ZN(n650) );
  NOR2_X1 U738 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n653), .A2(n652), .ZN(G290) );
  NAND2_X1 U740 ( .A1(G86), .A2(n654), .ZN(n656) );
  NAND2_X1 U741 ( .A1(G61), .A2(n668), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n657), .A2(G73), .ZN(n658) );
  XOR2_X1 U744 ( .A(KEYINPUT2), .B(n658), .Z(n659) );
  NOR2_X1 U745 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U746 ( .A1(G48), .A2(n663), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(G305) );
  NAND2_X1 U748 ( .A1(G651), .A2(G74), .ZN(n665) );
  NAND2_X1 U749 ( .A1(G49), .A2(n663), .ZN(n664) );
  NAND2_X1 U750 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U751 ( .A(KEYINPUT82), .B(n666), .ZN(n667) );
  NOR2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n669), .A2(G87), .ZN(n670) );
  NAND2_X1 U754 ( .A1(n671), .A2(n670), .ZN(G288) );
  XNOR2_X1 U755 ( .A(G166), .B(KEYINPUT19), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n987), .B(n679), .ZN(n674) );
  XOR2_X1 U757 ( .A(G305), .B(G288), .Z(n672) );
  XNOR2_X1 U758 ( .A(G290), .B(n672), .ZN(n673) );
  XNOR2_X1 U759 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U760 ( .A(n676), .B(n675), .ZN(n923) );
  XNOR2_X1 U761 ( .A(n677), .B(n923), .ZN(n678) );
  NAND2_X1 U762 ( .A1(n678), .A2(G868), .ZN(n681) );
  OR2_X1 U763 ( .A1(G868), .A2(n679), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U765 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U766 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U767 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U768 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XOR2_X1 U770 ( .A(KEYINPUT83), .B(G44), .Z(n686) );
  XNOR2_X1 U771 ( .A(KEYINPUT3), .B(n686), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U774 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U775 ( .A1(G96), .A2(n689), .ZN(n856) );
  NAND2_X1 U776 ( .A1(G2106), .A2(n856), .ZN(n693) );
  NAND2_X1 U777 ( .A1(G69), .A2(G120), .ZN(n690) );
  NOR2_X1 U778 ( .A1(G237), .A2(n690), .ZN(n691) );
  NAND2_X1 U779 ( .A1(G108), .A2(n691), .ZN(n857) );
  NAND2_X1 U780 ( .A1(G567), .A2(n857), .ZN(n692) );
  NAND2_X1 U781 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U782 ( .A(KEYINPUT84), .B(n694), .Z(G319) );
  INV_X1 U783 ( .A(G319), .ZN(n696) );
  NAND2_X1 U784 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n855) );
  NAND2_X1 U786 ( .A1(n855), .A2(G36), .ZN(G176) );
  INV_X1 U787 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT65), .ZN(n800) );
  NAND2_X1 U789 ( .A1(G160), .A2(G40), .ZN(n801) );
  NOR2_X1 U790 ( .A1(n800), .A2(n801), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G8), .A2(n733), .ZN(n748) );
  INV_X1 U792 ( .A(G8), .ZN(n751) );
  OR2_X1 U793 ( .A1(G1966), .A2(n751), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n707), .A2(n700), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n707), .A2(G2072), .ZN(n703) );
  INV_X1 U796 ( .A(G1956), .ZN(n1013) );
  NOR2_X1 U797 ( .A1(n752), .A2(n1013), .ZN(n704) );
  NOR2_X2 U798 ( .A1(n705), .A2(n704), .ZN(n721) );
  NOR2_X1 U799 ( .A1(n721), .A2(n987), .ZN(n706) );
  XNOR2_X1 U800 ( .A(n706), .B(KEYINPUT28), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n707), .A2(G2067), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n754), .A2(G1348), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n722) );
  NAND2_X1 U804 ( .A1(n722), .A2(n990), .ZN(n713) );
  XNOR2_X1 U805 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n710) );
  XNOR2_X1 U806 ( .A(n710), .B(KEYINPUT66), .ZN(n715) );
  NOR2_X1 U807 ( .A1(G1996), .A2(n715), .ZN(n711) );
  NOR2_X1 U808 ( .A1(n711), .A2(n1004), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n720) );
  INV_X1 U810 ( .A(G1341), .ZN(n1012) );
  NAND2_X1 U811 ( .A1(n1012), .A2(n715), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n714), .A2(n754), .ZN(n718) );
  INV_X1 U813 ( .A(G1996), .ZN(n967) );
  NOR2_X1 U814 ( .A1(n754), .A2(n967), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U816 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U817 ( .A1(n720), .A2(n719), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n721), .A2(n987), .ZN(n723) );
  NAND2_X1 U819 ( .A1(n723), .A2(n522), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n728), .B(KEYINPUT29), .ZN(n732) );
  INV_X1 U822 ( .A(G1961), .ZN(n1027) );
  NOR2_X1 U823 ( .A1(n752), .A2(n1027), .ZN(n730) );
  XNOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .ZN(n973) );
  NOR2_X1 U825 ( .A1(n754), .A2(n973), .ZN(n729) );
  NOR2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G171), .A2(n739), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n732), .A2(n731), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n746), .A2(n733), .ZN(n734) );
  NAND2_X1 U830 ( .A1(G8), .A2(n734), .ZN(n737) );
  XNOR2_X1 U831 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U832 ( .A1(G168), .A2(n738), .ZN(n741) );
  NOR2_X1 U833 ( .A1(G171), .A2(n739), .ZN(n740) );
  NOR2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U835 ( .A(KEYINPUT31), .B(n742), .Z(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n749) );
  INV_X1 U837 ( .A(n749), .ZN(n745) );
  NOR2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n767) );
  NAND2_X1 U840 ( .A1(G286), .A2(n749), .ZN(n750) );
  XNOR2_X1 U841 ( .A(n750), .B(KEYINPUT96), .ZN(n759) );
  OR2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n796) );
  NOR2_X1 U843 ( .A1(G1971), .A2(n796), .ZN(n753) );
  XNOR2_X1 U844 ( .A(KEYINPUT97), .B(n753), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n754), .A2(G2090), .ZN(n755) );
  NOR2_X1 U846 ( .A1(G166), .A2(n755), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n760), .A2(G8), .ZN(n761) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT32), .ZN(n769) );
  NAND2_X1 U851 ( .A1(n767), .A2(n769), .ZN(n764) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U853 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n765), .A2(n796), .ZN(n792) );
  NAND2_X1 U856 ( .A1(G288), .A2(G1976), .ZN(n766) );
  XOR2_X1 U857 ( .A(KEYINPUT98), .B(n766), .Z(n994) );
  NOR2_X1 U858 ( .A1(KEYINPUT99), .A2(n994), .ZN(n770) );
  AND2_X1 U859 ( .A1(n767), .A2(n770), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n784) );
  INV_X1 U861 ( .A(n770), .ZN(n772) );
  NOR2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n775) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U864 ( .A1(n775), .A2(n771), .ZN(n1002) );
  OR2_X1 U865 ( .A1(n772), .A2(n1002), .ZN(n782) );
  XOR2_X1 U866 ( .A(G1981), .B(G305), .Z(n998) );
  INV_X1 U867 ( .A(n998), .ZN(n780) );
  INV_X1 U868 ( .A(KEYINPUT99), .ZN(n774) );
  NAND2_X1 U869 ( .A1(n775), .A2(KEYINPUT33), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n775), .A2(KEYINPUT99), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n796), .A2(n778), .ZN(n779) );
  NOR2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n785) );
  AND2_X1 U875 ( .A1(n785), .A2(KEYINPUT33), .ZN(n788) );
  INV_X1 U876 ( .A(n788), .ZN(n781) );
  AND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n790) );
  INV_X1 U879 ( .A(n785), .ZN(n786) );
  NOR2_X1 U880 ( .A1(n796), .A2(n786), .ZN(n787) );
  OR2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U884 ( .A(KEYINPUT100), .B(n793), .ZN(n799) );
  NOR2_X1 U885 ( .A1(G1981), .A2(G305), .ZN(n794) );
  XOR2_X1 U886 ( .A(n794), .B(KEYINPUT24), .Z(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U888 ( .A(n797), .B(KEYINPUT92), .ZN(n798) );
  INV_X1 U889 ( .A(n801), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n800), .A2(n802), .ZN(n831) );
  NAND2_X1 U891 ( .A1(n907), .A2(G129), .ZN(n809) );
  NAND2_X1 U892 ( .A1(G117), .A2(n906), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G141), .A2(n902), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n903), .A2(G105), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT91), .B(n810), .Z(n899) );
  NAND2_X1 U900 ( .A1(G1996), .A2(n899), .ZN(n819) );
  NAND2_X1 U901 ( .A1(G119), .A2(n907), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G131), .A2(n902), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n906), .A2(G107), .ZN(n813) );
  XOR2_X1 U905 ( .A(KEYINPUT90), .B(n813), .Z(n814) );
  NOR2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n903), .A2(G95), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n913) );
  NAND2_X1 U909 ( .A1(G1991), .A2(n913), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n948) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n993) );
  NOR2_X1 U912 ( .A1(n948), .A2(n993), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n831), .A2(n820), .ZN(n833) );
  NAND2_X1 U914 ( .A1(G140), .A2(n902), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G104), .A2(n903), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U917 ( .A(KEYINPUT34), .B(n823), .ZN(n828) );
  NAND2_X1 U918 ( .A1(G116), .A2(n906), .ZN(n825) );
  NAND2_X1 U919 ( .A1(G128), .A2(n907), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U921 ( .A(n826), .B(KEYINPUT35), .Z(n827) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U923 ( .A(KEYINPUT36), .B(n829), .Z(n830) );
  XNOR2_X1 U924 ( .A(KEYINPUT89), .B(n830), .ZN(n917) );
  XNOR2_X1 U925 ( .A(G2067), .B(KEYINPUT37), .ZN(n843) );
  NOR2_X1 U926 ( .A1(n917), .A2(n843), .ZN(n947) );
  INV_X1 U927 ( .A(n831), .ZN(n845) );
  NAND2_X1 U928 ( .A1(n947), .A2(n845), .ZN(n842) );
  NAND2_X1 U929 ( .A1(n523), .A2(n834), .ZN(n849) );
  NOR2_X1 U930 ( .A1(G1996), .A2(n899), .ZN(n835) );
  XOR2_X1 U931 ( .A(KEYINPUT101), .B(n835), .Z(n952) );
  NOR2_X1 U932 ( .A1(G1986), .A2(G290), .ZN(n836) );
  NOR2_X1 U933 ( .A1(G1991), .A2(n913), .ZN(n944) );
  NOR2_X1 U934 ( .A1(n836), .A2(n944), .ZN(n837) );
  NOR2_X1 U935 ( .A1(n948), .A2(n837), .ZN(n838) );
  NOR2_X1 U936 ( .A1(n952), .A2(n838), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(KEYINPUT102), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(KEYINPUT39), .ZN(n841) );
  NAND2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n917), .A2(n843), .ZN(n949) );
  NAND2_X1 U941 ( .A1(n844), .A2(n949), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U943 ( .A(KEYINPUT103), .B(n847), .Z(n848) );
  NAND2_X1 U944 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U945 ( .A(n850), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U946 ( .A1(n851), .A2(G2106), .ZN(n852) );
  XOR2_X1 U947 ( .A(KEYINPUT105), .B(n852), .Z(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G661), .A2(n853), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G188) );
  XOR2_X1 U952 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U954 ( .A(G120), .ZN(G236) );
  INV_X1 U955 ( .A(G69), .ZN(G235) );
  NOR2_X1 U956 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U957 ( .A(G325), .ZN(G261) );
  XOR2_X1 U958 ( .A(KEYINPUT110), .B(G1986), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1981), .B(G1976), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n860), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U964 ( .A(G1971), .B(G1956), .Z(n864) );
  XNOR2_X1 U965 ( .A(G1966), .B(G1961), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U967 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U968 ( .A(KEYINPUT109), .B(G2474), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(G229) );
  XOR2_X1 U970 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n870) );
  XNOR2_X1 U971 ( .A(G2678), .B(KEYINPUT43), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U973 ( .A(KEYINPUT42), .B(G2072), .Z(n872) );
  XNOR2_X1 U974 ( .A(G2067), .B(G2090), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U977 ( .A(G2096), .B(G2100), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n878) );
  XOR2_X1 U979 ( .A(G2078), .B(G2084), .Z(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(G227) );
  NAND2_X1 U981 ( .A1(G124), .A2(n907), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n906), .A2(G112), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G136), .A2(n902), .ZN(n883) );
  NAND2_X1 U986 ( .A1(G100), .A2(n903), .ZN(n882) );
  NAND2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U988 ( .A1(n885), .A2(n884), .ZN(G162) );
  NAND2_X1 U989 ( .A1(n903), .A2(G106), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n886), .B(KEYINPUT112), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G142), .A2(n902), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n889), .B(KEYINPUT45), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G118), .A2(n906), .ZN(n891) );
  NAND2_X1 U995 ( .A1(G130), .A2(n907), .ZN(n890) );
  NAND2_X1 U996 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U997 ( .A(KEYINPUT111), .B(n892), .ZN(n893) );
  NAND2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U999 ( .A(n895), .B(G164), .ZN(n921) );
  XOR2_X1 U1000 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n897) );
  XNOR2_X1 U1001 ( .A(G162), .B(KEYINPUT114), .ZN(n896) );
  XNOR2_X1 U1002 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U1003 ( .A(KEYINPUT46), .B(n898), .ZN(n901) );
  XNOR2_X1 U1004 ( .A(n899), .B(KEYINPUT113), .ZN(n900) );
  XNOR2_X1 U1005 ( .A(n901), .B(n900), .ZN(n916) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n902), .ZN(n905) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n903), .ZN(n904) );
  NAND2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(G115), .A2(n906), .ZN(n909) );
  NAND2_X1 U1010 ( .A1(G127), .A2(n907), .ZN(n908) );
  NAND2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1012 ( .A(KEYINPUT47), .B(n910), .Z(n911) );
  NOR2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n936) );
  XNOR2_X1 U1014 ( .A(n936), .B(n913), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n914), .B(n941), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n917), .B(G160), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(n921), .B(n920), .Z(n922) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n922), .ZN(G395) );
  INV_X1 U1021 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U1022 ( .A(G286), .B(n923), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT116), .B(G301), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n924), .B(n990), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n926), .B(n925), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n927), .B(n1004), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(G37), .A2(n928), .ZN(G397) );
  NOR2_X1 U1028 ( .A1(G229), .A2(G227), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(n929), .B(KEYINPUT49), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(G401), .A2(n930), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n931), .A2(G319), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n932), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1035 ( .A(KEYINPUT118), .B(n935), .Z(G308) );
  INV_X1 U1036 ( .A(G308), .ZN(G225) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1038 ( .A(G164), .B(G2078), .ZN(n939) );
  XOR2_X1 U1039 ( .A(G2072), .B(n936), .Z(n937) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NAND2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n940), .B(KEYINPUT50), .ZN(n960) );
  XNOR2_X1 U1043 ( .A(G160), .B(G2084), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(KEYINPUT119), .B(n945), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n958) );
  INV_X1 U1048 ( .A(n948), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n953), .Z(n954) );
  XOR2_X1 U1053 ( .A(KEYINPUT120), .B(n954), .Z(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT52), .B(n961), .ZN(n962) );
  INV_X1 U1058 ( .A(KEYINPUT55), .ZN(n983) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n983), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n963), .A2(G29), .ZN(n1046) );
  XNOR2_X1 U1061 ( .A(G2084), .B(G34), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(n964), .B(KEYINPUT54), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(G35), .B(G2090), .ZN(n965) );
  NOR2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n981) );
  XNOR2_X1 U1065 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n979) );
  XOR2_X1 U1066 ( .A(G2072), .B(G33), .Z(n969) );
  XNOR2_X1 U1067 ( .A(n967), .B(G32), .ZN(n968) );
  NAND2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1069 ( .A(G26), .B(G2067), .ZN(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n977) );
  XOR2_X1 U1071 ( .A(G1991), .B(G25), .Z(n972) );
  NAND2_X1 U1072 ( .A1(n972), .A2(G28), .ZN(n975) );
  XOR2_X1 U1073 ( .A(G27), .B(n973), .Z(n974) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(n979), .B(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n983), .B(n982), .ZN(n985) );
  INV_X1 U1079 ( .A(G29), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n986), .ZN(n1044) );
  XNOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .ZN(n1010) );
  XNOR2_X1 U1083 ( .A(G1956), .B(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n988) );
  NAND2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(G1348), .B(n990), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1092 ( .A(KEYINPUT57), .B(n999), .Z(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G171), .B(G1961), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(n1012), .B(n1004), .Z(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1042) );
  INV_X1 U1100 ( .A(G16), .ZN(n1040) );
  XOR2_X1 U1101 ( .A(G1966), .B(G21), .Z(n1011) );
  XNOR2_X1 U1102 ( .A(KEYINPUT125), .B(n1011), .ZN(n1025) );
  XNOR2_X1 U1103 ( .A(n1012), .B(G19), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(n1013), .B(G20), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G6), .B(G1981), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(G4), .B(KEYINPUT123), .Z(n1019) );
  XNOR2_X1 U1109 ( .A(G1348), .B(KEYINPUT59), .ZN(n1018) );
  XNOR2_X1 U1110 ( .A(n1019), .B(n1018), .ZN(n1020) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1112 ( .A(KEYINPUT124), .B(n1022), .Z(n1023) );
  XOR2_X1 U1113 ( .A(KEYINPUT60), .B(n1023), .Z(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1115 ( .A(KEYINPUT126), .B(n1026), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(n1027), .B(G5), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(G1971), .B(G22), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(G24), .B(G1986), .ZN(n1030) );
  NOR2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  XOR2_X1 U1121 ( .A(G1976), .B(G23), .Z(n1032) );
  NAND2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1123 ( .A(KEYINPUT58), .B(n1034), .ZN(n1035) );
  NOR2_X1 U1124 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1125 ( .A(n1037), .B(KEYINPUT61), .Z(n1038) );
  XNOR2_X1 U1126 ( .A(KEYINPUT127), .B(n1038), .ZN(n1039) );
  NAND2_X1 U1127 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1128 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NOR2_X1 U1129 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1130 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XOR2_X1 U1131 ( .A(KEYINPUT62), .B(n1047), .Z(G311) );
  INV_X1 U1132 ( .A(G311), .ZN(G150) );
endmodule

