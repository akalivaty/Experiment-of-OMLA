

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(G2105), .ZN(n530) );
  NOR2_X2 U550 ( .A1(G164), .A2(G1384), .ZN(n755) );
  NOR2_X1 U551 ( .A1(n668), .A2(n667), .ZN(n685) );
  OR2_X1 U552 ( .A1(n673), .A2(n672), .ZN(n681) );
  BUF_X2 U553 ( .A(n980), .Z(n513) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n527), .Z(n980) );
  INV_X1 U555 ( .A(KEYINPUT28), .ZN(n686) );
  XNOR2_X1 U556 ( .A(n691), .B(n690), .ZN(n697) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n690) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XOR2_X1 U559 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U560 ( .A(KEYINPUT30), .B(KEYINPUT92), .ZN(n700) );
  XNOR2_X1 U561 ( .A(n701), .B(n700), .ZN(n702) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n706) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n628) );
  NOR2_X1 U564 ( .A1(G651), .A2(n621), .ZN(n627) );
  NOR2_X1 U565 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U566 ( .A(KEYINPUT71), .B(n526), .Z(G168) );
  XOR2_X1 U567 ( .A(G543), .B(KEYINPUT0), .Z(n621) );
  NAND2_X1 U568 ( .A1(G51), .A2(n627), .ZN(n516) );
  XNOR2_X1 U569 ( .A(KEYINPUT65), .B(G651), .ZN(n519) );
  NOR2_X1 U570 ( .A1(G543), .A2(n519), .ZN(n514) );
  XOR2_X2 U571 ( .A(KEYINPUT1), .B(n514), .Z(n631) );
  NAND2_X1 U572 ( .A1(G63), .A2(n631), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U574 ( .A(KEYINPUT6), .B(n517), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n628), .A2(G89), .ZN(n518) );
  XNOR2_X1 U576 ( .A(n518), .B(KEYINPUT4), .ZN(n521) );
  NOR2_X1 U577 ( .A1(n621), .A2(n519), .ZN(n635) );
  NAND2_X1 U578 ( .A1(G76), .A2(n635), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U580 ( .A(n522), .B(KEYINPUT5), .Z(n523) );
  XOR2_X1 U581 ( .A(KEYINPUT7), .B(n525), .Z(n526) );
  NAND2_X1 U582 ( .A1(G138), .A2(n513), .ZN(n529) );
  AND2_X4 U583 ( .A1(n530), .A2(G2104), .ZN(n978) );
  NAND2_X1 U584 ( .A1(G102), .A2(n978), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n534) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n975) );
  NAND2_X1 U587 ( .A1(G114), .A2(n975), .ZN(n532) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n530), .ZN(n976) );
  NAND2_X1 U589 ( .A1(G126), .A2(n976), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U592 ( .A1(G101), .A2(n978), .ZN(n535) );
  XNOR2_X1 U593 ( .A(n535), .B(KEYINPUT64), .ZN(n537) );
  INV_X1 U594 ( .A(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U595 ( .A(n537), .B(n536), .ZN(n539) );
  NAND2_X1 U596 ( .A1(G137), .A2(n513), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U598 ( .A1(G113), .A2(n975), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G125), .A2(n976), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X2 U601 ( .A1(n543), .A2(n542), .ZN(G160) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  NAND2_X1 U605 ( .A1(G53), .A2(n627), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G65), .A2(n631), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n628), .A2(G91), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G78), .A2(n635), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n684) );
  INV_X1 U612 ( .A(n684), .ZN(G299) );
  XNOR2_X1 U613 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n628), .A2(G90), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G77), .A2(n635), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT9), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G52), .A2(n627), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G64), .A2(n631), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n558), .A2(n557), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n559) );
  XOR2_X1 U625 ( .A(n559), .B(KEYINPUT10), .Z(n1017) );
  NAND2_X1 U626 ( .A1(n1017), .A2(G567), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  XOR2_X1 U628 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n562) );
  NAND2_X1 U629 ( .A1(G56), .A2(n631), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n628), .A2(G81), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G68), .A2(n635), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n627), .A2(G43), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n916) );
  INV_X1 U639 ( .A(G860), .ZN(n582) );
  OR2_X1 U640 ( .A1(n916), .A2(n582), .ZN(G153) );
  NAND2_X1 U641 ( .A1(G868), .A2(G301), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n628), .A2(G92), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G66), .A2(n631), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n627), .A2(G54), .ZN(n574) );
  NAND2_X1 U646 ( .A1(G79), .A2(n635), .ZN(n573) );
  NAND2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U649 ( .A(KEYINPUT15), .B(n577), .ZN(n972) );
  INV_X1 U650 ( .A(G868), .ZN(n648) );
  NAND2_X1 U651 ( .A1(n972), .A2(n648), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(G284) );
  NOR2_X1 U653 ( .A1(G286), .A2(n648), .ZN(n581) );
  NOR2_X1 U654 ( .A1(G868), .A2(G299), .ZN(n580) );
  NOR2_X1 U655 ( .A1(n581), .A2(n580), .ZN(G297) );
  NAND2_X1 U656 ( .A1(n582), .A2(G559), .ZN(n583) );
  INV_X1 U657 ( .A(n972), .ZN(n673) );
  NAND2_X1 U658 ( .A1(n583), .A2(n673), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U660 ( .A1(n972), .A2(n648), .ZN(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT72), .B(n585), .Z(n586) );
  NOR2_X1 U662 ( .A1(G559), .A2(n586), .ZN(n588) );
  NOR2_X1 U663 ( .A1(G868), .A2(n916), .ZN(n587) );
  NOR2_X1 U664 ( .A1(n588), .A2(n587), .ZN(G282) );
  NAND2_X1 U665 ( .A1(G123), .A2(n976), .ZN(n589) );
  XOR2_X1 U666 ( .A(KEYINPUT18), .B(n589), .Z(n590) );
  XNOR2_X1 U667 ( .A(n590), .B(KEYINPUT73), .ZN(n592) );
  NAND2_X1 U668 ( .A1(G111), .A2(n975), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G135), .A2(n513), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G99), .A2(n978), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n989) );
  XNOR2_X1 U674 ( .A(n989), .B(G2096), .ZN(n597) );
  INV_X1 U675 ( .A(G2100), .ZN(n937) );
  NAND2_X1 U676 ( .A1(n597), .A2(n937), .ZN(G156) );
  NAND2_X1 U677 ( .A1(n673), .A2(G559), .ZN(n645) );
  XNOR2_X1 U678 ( .A(n916), .B(n645), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n598), .A2(G860), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n628), .A2(G93), .ZN(n600) );
  NAND2_X1 U681 ( .A1(G67), .A2(n631), .ZN(n599) );
  NAND2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n627), .A2(G55), .ZN(n602) );
  NAND2_X1 U684 ( .A1(G80), .A2(n635), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  OR2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n647) );
  XOR2_X1 U687 ( .A(n605), .B(n647), .Z(G145) );
  NAND2_X1 U688 ( .A1(G48), .A2(n627), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G86), .A2(n628), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n635), .A2(G73), .ZN(n608) );
  XOR2_X1 U692 ( .A(KEYINPUT2), .B(n608), .Z(n609) );
  NOR2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G61), .A2(n631), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(G305) );
  NAND2_X1 U696 ( .A1(G62), .A2(n631), .ZN(n613) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT74), .ZN(n615) );
  NAND2_X1 U698 ( .A1(G50), .A2(n627), .ZN(n614) );
  NAND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U700 ( .A(KEYINPUT75), .B(n616), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n635), .A2(G75), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n628), .A2(G88), .ZN(n617) );
  AND2_X1 U703 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(G303) );
  NAND2_X1 U705 ( .A1(G87), .A2(n621), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n631), .A2(n624), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(G49), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G47), .A2(n627), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G85), .A2(n628), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n631), .A2(G60), .ZN(n632) );
  XOR2_X1 U715 ( .A(KEYINPUT66), .B(n632), .Z(n633) );
  NOR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G72), .A2(n635), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(G290) );
  XOR2_X1 U719 ( .A(n647), .B(G305), .Z(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT19), .B(n684), .Z(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(G288), .ZN(n639) );
  XOR2_X1 U722 ( .A(G303), .B(n639), .Z(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(G290), .ZN(n641) );
  XNOR2_X1 U724 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(n916), .ZN(n970) );
  XOR2_X1 U726 ( .A(n970), .B(KEYINPUT76), .Z(n644) );
  XNOR2_X1 U727 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n646), .A2(G868), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n651), .Z(n652) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n652), .ZN(n653) );
  XNOR2_X1 U734 ( .A(KEYINPUT21), .B(n653), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n654), .A2(G2072), .ZN(n655) );
  XOR2_X1 U736 ( .A(KEYINPUT77), .B(n655), .Z(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U738 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NAND2_X1 U739 ( .A1(G661), .A2(G483), .ZN(n663) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT22), .B(n656), .Z(n657) );
  NOR2_X1 U742 ( .A1(G218), .A2(n657), .ZN(n658) );
  NAND2_X1 U743 ( .A1(G96), .A2(n658), .ZN(n935) );
  NAND2_X1 U744 ( .A1(n935), .A2(G2106), .ZN(n662) );
  NAND2_X1 U745 ( .A1(G69), .A2(G120), .ZN(n659) );
  NOR2_X1 U746 ( .A1(G237), .A2(n659), .ZN(n660) );
  NAND2_X1 U747 ( .A1(G108), .A2(n660), .ZN(n934) );
  NAND2_X1 U748 ( .A1(n934), .A2(G567), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n662), .A2(n661), .ZN(n1016) );
  NOR2_X1 U750 ( .A1(n663), .A2(n1016), .ZN(n664) );
  XNOR2_X1 U751 ( .A(n664), .B(KEYINPUT78), .ZN(n812) );
  NAND2_X1 U752 ( .A1(G36), .A2(n812), .ZN(G176) );
  INV_X1 U753 ( .A(G303), .ZN(G166) );
  NAND2_X1 U754 ( .A1(G160), .A2(G40), .ZN(n754) );
  INV_X1 U755 ( .A(n754), .ZN(n665) );
  NAND2_X2 U756 ( .A1(n755), .A2(n665), .ZN(n711) );
  XNOR2_X2 U757 ( .A(n711), .B(KEYINPUT89), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n692), .A2(G2072), .ZN(n666) );
  XNOR2_X1 U759 ( .A(n666), .B(KEYINPUT27), .ZN(n668) );
  INV_X1 U760 ( .A(G1956), .ZN(n954) );
  NOR2_X1 U761 ( .A1(n954), .A2(n692), .ZN(n667) );
  NAND2_X1 U762 ( .A1(n685), .A2(n684), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G2067), .A2(n692), .ZN(n669) );
  XNOR2_X1 U764 ( .A(n669), .B(KEYINPUT91), .ZN(n671) );
  AND2_X1 U765 ( .A1(G1348), .A2(n711), .ZN(n670) );
  NOR2_X1 U766 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U767 ( .A1(n673), .A2(n672), .ZN(n679) );
  INV_X1 U768 ( .A(G1996), .ZN(n949) );
  NOR2_X1 U769 ( .A1(n711), .A2(n949), .ZN(n674) );
  XOR2_X1 U770 ( .A(n674), .B(KEYINPUT26), .Z(n676) );
  NAND2_X1 U771 ( .A1(n711), .A2(G1341), .ZN(n675) );
  NAND2_X1 U772 ( .A1(n676), .A2(n675), .ZN(n677) );
  OR2_X1 U773 ( .A1(n916), .A2(n677), .ZN(n678) );
  NAND2_X1 U774 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U775 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U776 ( .A1(n683), .A2(n682), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U780 ( .A(G1961), .ZN(n946) );
  NAND2_X1 U781 ( .A1(n946), .A2(n711), .ZN(n694) );
  XNOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .ZN(n831) );
  NAND2_X1 U783 ( .A1(n692), .A2(n831), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n703) );
  AND2_X1 U785 ( .A1(n703), .A2(G171), .ZN(n695) );
  XOR2_X1 U786 ( .A(KEYINPUT90), .B(n695), .Z(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n709) );
  NAND2_X1 U788 ( .A1(G8), .A2(n711), .ZN(n747) );
  NOR2_X1 U789 ( .A1(G1966), .A2(n747), .ZN(n723) );
  NOR2_X1 U790 ( .A1(n711), .A2(G2084), .ZN(n698) );
  XNOR2_X1 U791 ( .A(n698), .B(KEYINPUT88), .ZN(n720) );
  NOR2_X1 U792 ( .A1(n723), .A2(n720), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n699), .A2(G8), .ZN(n701) );
  NOR2_X1 U794 ( .A1(G168), .A2(n702), .ZN(n705) );
  NOR2_X1 U795 ( .A1(G171), .A2(n703), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n721) );
  NAND2_X1 U799 ( .A1(n721), .A2(G286), .ZN(n718) );
  INV_X1 U800 ( .A(G8), .ZN(n716) );
  NOR2_X1 U801 ( .A1(G1971), .A2(n747), .ZN(n710) );
  XNOR2_X1 U802 ( .A(KEYINPUT93), .B(n710), .ZN(n714) );
  NOR2_X1 U803 ( .A1(G2090), .A2(n711), .ZN(n712) );
  NOR2_X1 U804 ( .A1(G166), .A2(n712), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U808 ( .A(n719), .B(KEYINPUT32), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n720), .A2(G8), .ZN(n725) );
  INV_X1 U810 ( .A(n721), .ZN(n722) );
  NOR2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n743) );
  NOR2_X1 U814 ( .A1(G1976), .A2(G288), .ZN(n909) );
  INV_X1 U815 ( .A(n909), .ZN(n730) );
  NOR2_X1 U816 ( .A1(G1971), .A2(G303), .ZN(n728) );
  XOR2_X1 U817 ( .A(n728), .B(KEYINPUT94), .Z(n729) );
  AND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U819 ( .A1(n743), .A2(n731), .ZN(n732) );
  XNOR2_X1 U820 ( .A(n732), .B(KEYINPUT95), .ZN(n733) );
  NAND2_X1 U821 ( .A1(G1976), .A2(G288), .ZN(n910) );
  NAND2_X1 U822 ( .A1(n733), .A2(n910), .ZN(n734) );
  XNOR2_X1 U823 ( .A(KEYINPUT96), .B(n734), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n735), .A2(n747), .ZN(n736) );
  NOR2_X1 U825 ( .A1(KEYINPUT33), .A2(n736), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n909), .A2(KEYINPUT33), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n747), .A2(n737), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U829 ( .A(G1981), .B(G305), .Z(n921) );
  NAND2_X1 U830 ( .A1(n740), .A2(n921), .ZN(n751) );
  NOR2_X1 U831 ( .A1(G2090), .A2(G303), .ZN(n741) );
  NAND2_X1 U832 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U834 ( .A1(n747), .A2(n744), .ZN(n749) );
  NOR2_X1 U835 ( .A1(G1981), .A2(G305), .ZN(n745) );
  XOR2_X1 U836 ( .A(n745), .B(KEYINPUT24), .Z(n746) );
  NOR2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n753) );
  INV_X1 U840 ( .A(KEYINPUT97), .ZN(n752) );
  XNOR2_X1 U841 ( .A(n753), .B(n752), .ZN(n792) );
  XNOR2_X1 U842 ( .A(G1986), .B(G290), .ZN(n913) );
  NOR2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n804) );
  NAND2_X1 U844 ( .A1(n913), .A2(n804), .ZN(n756) );
  XOR2_X1 U845 ( .A(n756), .B(KEYINPUT79), .Z(n790) );
  NAND2_X1 U846 ( .A1(n978), .A2(G105), .ZN(n758) );
  XNOR2_X1 U847 ( .A(KEYINPUT38), .B(KEYINPUT86), .ZN(n757) );
  XNOR2_X1 U848 ( .A(n758), .B(n757), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G117), .A2(n975), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G129), .A2(n976), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n763) );
  NAND2_X1 U852 ( .A1(G141), .A2(n513), .ZN(n761) );
  XNOR2_X1 U853 ( .A(KEYINPUT87), .B(n761), .ZN(n762) );
  NOR2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n999) );
  NAND2_X1 U856 ( .A1(G1996), .A2(n999), .ZN(n774) );
  XOR2_X1 U857 ( .A(G1991), .B(KEYINPUT85), .Z(n826) );
  NAND2_X1 U858 ( .A1(G119), .A2(n976), .ZN(n767) );
  NAND2_X1 U859 ( .A1(G131), .A2(n513), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n975), .A2(G107), .ZN(n768) );
  XOR2_X1 U862 ( .A(KEYINPUT84), .B(n768), .Z(n769) );
  NOR2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n978), .A2(G95), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n992) );
  NAND2_X1 U866 ( .A1(n826), .A2(n992), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n884) );
  NAND2_X1 U868 ( .A1(n884), .A2(n804), .ZN(n788) );
  NAND2_X1 U869 ( .A1(n513), .A2(G140), .ZN(n775) );
  XNOR2_X1 U870 ( .A(n775), .B(KEYINPUT80), .ZN(n777) );
  NAND2_X1 U871 ( .A1(G104), .A2(n978), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U873 ( .A(KEYINPUT34), .B(n778), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n976), .A2(G128), .ZN(n779) );
  XNOR2_X1 U875 ( .A(KEYINPUT81), .B(n779), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n975), .A2(G116), .ZN(n780) );
  XOR2_X1 U877 ( .A(KEYINPUT82), .B(n780), .Z(n781) );
  NOR2_X1 U878 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U879 ( .A(n783), .B(KEYINPUT35), .ZN(n784) );
  NOR2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n787) );
  XOR2_X1 U881 ( .A(KEYINPUT83), .B(KEYINPUT36), .Z(n786) );
  XOR2_X1 U882 ( .A(n787), .B(n786), .Z(n993) );
  XOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .Z(n803) );
  AND2_X1 U884 ( .A1(n993), .A2(n803), .ZN(n888) );
  NAND2_X1 U885 ( .A1(n888), .A2(n804), .ZN(n793) );
  AND2_X1 U886 ( .A1(n788), .A2(n793), .ZN(n789) );
  AND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n808) );
  INV_X1 U889 ( .A(n793), .ZN(n802) );
  NOR2_X1 U890 ( .A1(n999), .A2(G1996), .ZN(n794) );
  XNOR2_X1 U891 ( .A(n794), .B(KEYINPUT98), .ZN(n880) );
  NOR2_X1 U892 ( .A1(n826), .A2(n992), .ZN(n882) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n795) );
  XOR2_X1 U894 ( .A(n795), .B(KEYINPUT99), .Z(n796) );
  NOR2_X1 U895 ( .A1(n882), .A2(n796), .ZN(n797) );
  NOR2_X1 U896 ( .A1(n884), .A2(n797), .ZN(n798) );
  NOR2_X1 U897 ( .A1(n880), .A2(n798), .ZN(n799) );
  XNOR2_X1 U898 ( .A(KEYINPUT39), .B(n799), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n800), .A2(n804), .ZN(n801) );
  OR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n993), .A2(n803), .ZN(n893) );
  NAND2_X1 U902 ( .A1(n893), .A2(n804), .ZN(n805) );
  AND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U905 ( .A(n809), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n1017), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n810) );
  NAND2_X1 U908 ( .A1(G661), .A2(n810), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n811) );
  NAND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(G188) );
  XOR2_X1 U911 ( .A(G96), .B(KEYINPUT102), .Z(G221) );
  NAND2_X1 U913 ( .A1(G100), .A2(n978), .ZN(n813) );
  XNOR2_X1 U914 ( .A(n813), .B(KEYINPUT106), .ZN(n816) );
  NAND2_X1 U915 ( .A1(G136), .A2(n513), .ZN(n814) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(n814), .Z(n815) );
  NAND2_X1 U917 ( .A1(n816), .A2(n815), .ZN(n821) );
  NAND2_X1 U918 ( .A1(G124), .A2(n976), .ZN(n817) );
  XNOR2_X1 U919 ( .A(n817), .B(KEYINPUT44), .ZN(n819) );
  NAND2_X1 U920 ( .A1(n975), .A2(G112), .ZN(n818) );
  NAND2_X1 U921 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U922 ( .A1(n821), .A2(n820), .ZN(G162) );
  XOR2_X1 U923 ( .A(KEYINPUT121), .B(n949), .Z(n822) );
  XNOR2_X1 U924 ( .A(n822), .B(G32), .ZN(n830) );
  XNOR2_X1 U925 ( .A(G2067), .B(G26), .ZN(n824) );
  XNOR2_X1 U926 ( .A(G33), .B(G2072), .ZN(n823) );
  NOR2_X1 U927 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U928 ( .A1(G28), .A2(n825), .ZN(n828) );
  XNOR2_X1 U929 ( .A(G25), .B(n826), .ZN(n827) );
  NOR2_X1 U930 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U931 ( .A1(n830), .A2(n829), .ZN(n833) );
  XOR2_X1 U932 ( .A(G27), .B(n831), .Z(n832) );
  NOR2_X1 U933 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U934 ( .A(KEYINPUT53), .B(n834), .Z(n837) );
  XOR2_X1 U935 ( .A(G34), .B(KEYINPUT54), .Z(n835) );
  XNOR2_X1 U936 ( .A(G2084), .B(n835), .ZN(n836) );
  NAND2_X1 U937 ( .A1(n837), .A2(n836), .ZN(n839) );
  XNOR2_X1 U938 ( .A(G35), .B(G2090), .ZN(n838) );
  NOR2_X1 U939 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT55), .B(n840), .Z(n842) );
  INV_X1 U941 ( .A(G29), .ZN(n900) );
  XOR2_X1 U942 ( .A(n900), .B(KEYINPUT122), .Z(n841) );
  NOR2_X1 U943 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U944 ( .A(KEYINPUT123), .B(n843), .ZN(n905) );
  XOR2_X1 U945 ( .A(G5), .B(G1961), .Z(n856) );
  XNOR2_X1 U946 ( .A(G1348), .B(KEYINPUT59), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n844), .B(G4), .ZN(n848) );
  XNOR2_X1 U948 ( .A(G1341), .B(G19), .ZN(n846) );
  XNOR2_X1 U949 ( .A(G1981), .B(G6), .ZN(n845) );
  NOR2_X1 U950 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n851) );
  XNOR2_X1 U952 ( .A(G20), .B(G1956), .ZN(n849) );
  XNOR2_X1 U953 ( .A(KEYINPUT126), .B(n849), .ZN(n850) );
  NOR2_X1 U954 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(KEYINPUT60), .B(n852), .Z(n854) );
  XNOR2_X1 U956 ( .A(G1966), .B(G21), .ZN(n853) );
  NOR2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n863) );
  XNOR2_X1 U959 ( .A(G1971), .B(G22), .ZN(n858) );
  XNOR2_X1 U960 ( .A(G23), .B(G1976), .ZN(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n860) );
  XOR2_X1 U962 ( .A(G1986), .B(G24), .Z(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U964 ( .A(KEYINPUT58), .B(n861), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U966 ( .A(KEYINPUT61), .B(n864), .ZN(n865) );
  INV_X1 U967 ( .A(G16), .ZN(n906) );
  NAND2_X1 U968 ( .A1(n865), .A2(n906), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n866), .A2(G11), .ZN(n903) );
  NAND2_X1 U970 ( .A1(G115), .A2(n975), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G127), .A2(n976), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n869), .B(KEYINPUT47), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G103), .A2(n978), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G139), .A2(n513), .ZN(n872) );
  XNOR2_X1 U977 ( .A(KEYINPUT111), .B(n872), .ZN(n873) );
  NOR2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n991) );
  XNOR2_X1 U979 ( .A(G2072), .B(n991), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n875), .B(KEYINPUT119), .ZN(n877) );
  XOR2_X1 U981 ( .A(G2078), .B(G164), .Z(n876) );
  NOR2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U983 ( .A(KEYINPUT50), .B(n878), .Z(n896) );
  XOR2_X1 U984 ( .A(G2090), .B(G162), .Z(n879) );
  NOR2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U986 ( .A(KEYINPUT51), .B(n881), .Z(n891) );
  NOR2_X1 U987 ( .A1(n882), .A2(n989), .ZN(n886) );
  XOR2_X1 U988 ( .A(G160), .B(G2084), .Z(n883) );
  NOR2_X1 U989 ( .A1(n884), .A2(n883), .ZN(n885) );
  NAND2_X1 U990 ( .A1(n886), .A2(n885), .ZN(n887) );
  NOR2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U992 ( .A(KEYINPUT117), .B(n889), .Z(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT118), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(n897), .B(KEYINPUT52), .Z(n898) );
  XNOR2_X1 U998 ( .A(KEYINPUT120), .B(n898), .ZN(n899) );
  NOR2_X1 U999 ( .A1(KEYINPUT55), .A2(n899), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n932) );
  XNOR2_X1 U1003 ( .A(n906), .B(KEYINPUT56), .ZN(n930) );
  XOR2_X1 U1004 ( .A(G301), .B(G1961), .Z(n920) );
  XOR2_X1 U1005 ( .A(G1348), .B(n972), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(KEYINPUT124), .ZN(n915) );
  XOR2_X1 U1007 ( .A(G299), .B(n954), .Z(n908) );
  NOR2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(G1341), .B(n916), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n927) );
  XOR2_X1 U1015 ( .A(G303), .B(G1971), .Z(n925) );
  XNOR2_X1 U1016 ( .A(G1966), .B(G168), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(n923), .B(KEYINPUT57), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1021 ( .A(KEYINPUT125), .B(n928), .Z(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(n933), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1025 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1026 ( .A(G120), .ZN(G236) );
  INV_X1 U1027 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1029 ( .A(n936), .B(KEYINPUT103), .Z(G325) );
  INV_X1 U1030 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1031 ( .A(n937), .B(G2096), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G2072), .B(G2090), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n939), .B(n938), .ZN(n943) );
  XOR2_X1 U1034 ( .A(G2678), .B(KEYINPUT42), .Z(n941) );
  XNOR2_X1 U1035 ( .A(G2067), .B(KEYINPUT43), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n941), .B(n940), .ZN(n942) );
  XOR2_X1 U1037 ( .A(n943), .B(n942), .Z(n945) );
  XNOR2_X1 U1038 ( .A(G2078), .B(G2084), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n945), .B(n944), .ZN(G227) );
  XOR2_X1 U1040 ( .A(G1986), .B(n946), .Z(n958) );
  XOR2_X1 U1041 ( .A(G2474), .B(G1976), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G1971), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n953) );
  XOR2_X1 U1044 ( .A(KEYINPUT104), .B(G1981), .Z(n951) );
  XOR2_X1 U1045 ( .A(n949), .B(G1991), .Z(n950) );
  XNOR2_X1 U1046 ( .A(n951), .B(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(n953), .B(n952), .Z(n956) );
  XOR2_X1 U1048 ( .A(n954), .B(KEYINPUT41), .Z(n955) );
  XNOR2_X1 U1049 ( .A(n956), .B(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n958), .B(n957), .ZN(G229) );
  XNOR2_X1 U1051 ( .A(G2443), .B(G1341), .ZN(n967) );
  XNOR2_X1 U1052 ( .A(G2430), .B(G2435), .ZN(n965) );
  XOR2_X1 U1053 ( .A(KEYINPUT100), .B(G2454), .Z(n960) );
  XNOR2_X1 U1054 ( .A(G2427), .B(G2451), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n960), .B(n959), .ZN(n961) );
  XOR2_X1 U1056 ( .A(n961), .B(G2446), .Z(n963) );
  XNOR2_X1 U1057 ( .A(G1348), .B(G2438), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(n963), .B(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n965), .B(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n967), .B(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n968), .A2(G14), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT101), .B(n969), .ZN(G401) );
  XOR2_X1 U1063 ( .A(G301), .B(G286), .Z(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(n970), .ZN(n973) );
  XOR2_X1 U1065 ( .A(n973), .B(n972), .Z(n974) );
  NOR2_X1 U1066 ( .A1(G37), .A2(n974), .ZN(G397) );
  NAND2_X1 U1067 ( .A1(G118), .A2(n975), .ZN(n988) );
  NAND2_X1 U1068 ( .A1(n976), .A2(G130), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(KEYINPUT107), .B(n977), .ZN(n986) );
  NAND2_X1 U1070 ( .A1(n978), .A2(G106), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT108), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(G142), .A2(n513), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(KEYINPUT109), .B(n983), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT45), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n990), .B(n989), .ZN(n997) );
  XNOR2_X1 U1079 ( .A(n992), .B(n991), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(n993), .B(G160), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(n995), .B(n994), .ZN(n996) );
  XOR2_X1 U1082 ( .A(n997), .B(n996), .Z(n998) );
  XNOR2_X1 U1083 ( .A(n999), .B(n998), .ZN(n1004) );
  XOR2_X1 U1084 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n1001) );
  XNOR2_X1 U1085 ( .A(G162), .B(KEYINPUT48), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G164), .B(n1002), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(n1004), .B(n1003), .ZN(n1005) );
  NOR2_X1 U1089 ( .A1(G37), .A2(n1005), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(KEYINPUT112), .B(n1006), .ZN(G395) );
  XNOR2_X1 U1091 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n1008) );
  NOR2_X1 U1092 ( .A1(G227), .A2(G229), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT114), .B(n1009), .Z(n1012) );
  NOR2_X1 U1095 ( .A1(G401), .A2(n1016), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(KEYINPUT113), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(KEYINPUT116), .B(n1013), .ZN(n1015) );
  NOR2_X1 U1099 ( .A1(G397), .A2(G395), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(G225) );
  INV_X1 U1101 ( .A(G225), .ZN(G308) );
  INV_X1 U1102 ( .A(n1016), .ZN(G319) );
  INV_X1 U1103 ( .A(G108), .ZN(G238) );
  INV_X1 U1104 ( .A(n1017), .ZN(G223) );
endmodule

