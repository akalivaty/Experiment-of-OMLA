//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT80), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT79), .Z(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT27), .B(G183gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT69), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT28), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT68), .B(G183gat), .Z(new_n224));
  AOI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(KEYINPUT27), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n225), .B2(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n217), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  INV_X1    g027(.A(new_n213), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(KEYINPUT23), .B2(new_n214), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT65), .B1(new_n211), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n214), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n230), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(KEYINPUT64), .A3(new_n241), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n236), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n230), .B1(new_n233), .B2(new_n235), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n228), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n233), .A2(new_n235), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n213), .B(KEYINPUT67), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT25), .B1(new_n211), .B2(new_n232), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n240), .B1(new_n224), .B2(G190gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n227), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n207), .B1(new_n256), .B2(KEYINPUT29), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT78), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT77), .B(G218gat), .ZN(new_n260));
  INV_X1    g059(.A(G211gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n262), .B2(new_n263), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n263), .ZN(new_n269));
  INV_X1    g068(.A(new_n264), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT78), .A3(new_n265), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n207), .ZN(new_n275));
  INV_X1    g074(.A(new_n255), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n236), .A3(new_n244), .A4(new_n245), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(new_n228), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n275), .B1(new_n279), .B2(new_n227), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n257), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n257), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n205), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n257), .A2(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n273), .ZN(new_n285));
  INV_X1    g084(.A(new_n205), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n257), .A2(new_n274), .A3(new_n280), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n288), .A3(KEYINPUT30), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n285), .A2(new_n290), .A3(new_n287), .A4(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT82), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  INV_X1    g094(.A(G148gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT2), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G155gat), .B(G162gat), .Z(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n302), .C1(new_n303), .C2(KEYINPUT81), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n297), .A3(new_n298), .ZN(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n297), .A2(KEYINPUT81), .A3(new_n298), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G113gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n310), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G127gat), .B(G134gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT70), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n311), .A2(G120gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n325));
  NAND2_X1  g124(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n316), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n321), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n309), .A2(new_n324), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n323), .B1(new_n327), .B2(new_n331), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(new_n309), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n294), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n335), .B2(new_n309), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n309), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n332), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n304), .A2(new_n308), .A3(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n294), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(KEYINPUT5), .B(new_n337), .C1(new_n341), .C2(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n338), .A2(KEYINPUT83), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n339), .A3(new_n309), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n351), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G1gat), .B(G29gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n349), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n349), .A2(new_n357), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n361), .B(KEYINPUT87), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n349), .A2(new_n357), .A3(new_n369), .A4(new_n361), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n363), .A2(new_n367), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n361), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(KEYINPUT6), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n292), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT90), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT35), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n379));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n343), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n273), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n309), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n271), .B2(new_n265), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n342), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT85), .B(KEYINPUT29), .C1(new_n271), .C2(new_n265), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n382), .A2(new_n268), .A3(new_n272), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n384), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n383), .A2(new_n389), .B1(new_n392), .B2(new_n380), .ZN(new_n393));
  INV_X1    g192(.A(G22gat), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n379), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT31), .B(G50gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n389), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n392), .A2(new_n380), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n400), .A2(new_n401), .A3(new_n394), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n395), .A2(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G22gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n393), .A2(new_n394), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(new_n379), .A3(new_n407), .A4(new_n398), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n256), .A2(new_n344), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n335), .B1(new_n279), .B2(new_n227), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G15gat), .B(G43gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT73), .ZN(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT74), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n424), .B2(new_n422), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(KEYINPUT32), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n414), .B1(new_n410), .B2(new_n411), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT34), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT34), .B(new_n414), .C1(new_n410), .C2(new_n411), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n423), .A3(new_n427), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n378), .A2(new_n409), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n292), .A2(KEYINPUT90), .A3(new_n374), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n377), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n428), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n423), .A2(KEYINPUT75), .A3(new_n427), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n433), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n364), .A2(new_n372), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n363), .A2(new_n445), .A3(new_n368), .A4(new_n370), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n289), .A2(new_n291), .B1(new_n373), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n444), .A2(new_n447), .A3(new_n436), .A4(new_n409), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n439), .A2(new_n440), .B1(new_n448), .B2(KEYINPUT35), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n377), .A2(new_n437), .A3(KEYINPUT91), .A4(new_n438), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n355), .A2(new_n351), .A3(new_n346), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n294), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n365), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT89), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n456), .A3(new_n365), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n294), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT39), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n334), .A2(new_n336), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(new_n347), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n367), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n455), .A2(new_n457), .B1(new_n459), .B2(new_n462), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n289), .B(new_n291), .C1(new_n467), .C2(KEYINPUT40), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT37), .B1(new_n281), .B2(new_n282), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n285), .A2(new_n471), .A3(new_n287), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n472), .A3(new_n205), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n288), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n371), .A2(new_n373), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n470), .A2(new_n472), .A3(new_n474), .A4(new_n205), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n409), .B1(new_n469), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n409), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n447), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n436), .A2(KEYINPUT36), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT76), .B1(new_n444), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n434), .A2(new_n436), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n444), .A2(new_n484), .A3(KEYINPUT76), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n449), .A2(new_n450), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT104), .ZN(new_n493));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(KEYINPUT12), .Z(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n500), .A2(G1gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT16), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n502), .B2(G1gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G8gat), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  OR3_X1    g311(.A1(KEYINPUT93), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT14), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(KEYINPUT93), .C1(G29gat), .C2(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n518), .B(new_n519), .C1(new_n510), .C2(KEYINPUT15), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n512), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G43gat), .ZN(new_n523));
  INV_X1    g322(.A(G43gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G50gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n526), .A2(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(new_n511), .A3(new_n515), .A4(new_n518), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n521), .A2(new_n529), .A3(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n509), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n508), .A2(new_n530), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT95), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n535), .B(KEYINPUT13), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT96), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n505), .A2(new_n521), .A3(new_n529), .A4(new_n507), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n508), .A2(KEYINPUT96), .A3(new_n530), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n542), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n499), .B1(new_n539), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n549), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n552), .A2(new_n543), .B1(new_n540), .B2(new_n541), .ZN(new_n553));
  INV_X1    g352(.A(new_n499), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n537), .A2(KEYINPUT95), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n537), .A2(KEYINPUT95), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  AND4_X1   g368(.A1(new_n562), .A2(new_n565), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n560), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n562), .A2(new_n565), .A3(new_n568), .A4(new_n569), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT99), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n573), .A2(KEYINPUT100), .A3(new_n574), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT100), .B1(new_n573), .B2(new_n574), .ZN(new_n577));
  OAI22_X1  g376(.A1(new_n572), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT101), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n570), .A2(new_n560), .A3(new_n571), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT99), .B1(new_n573), .B2(new_n574), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(new_n577), .C2(new_n576), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n533), .A3(new_n532), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n530), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G190gat), .B(G218gat), .Z(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n591), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G57gat), .B(G64gat), .Z(new_n596));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n597), .B1(new_n596), .B2(new_n601), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n605));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n602), .B2(new_n603), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n596), .A2(new_n601), .ZN(new_n610));
  INV_X1    g409(.A(new_n597), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT98), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n508), .B1(new_n615), .B2(KEYINPUT21), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n607), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT97), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n595), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n578), .B1(new_n603), .B2(new_n602), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n570), .A2(KEYINPUT102), .A3(new_n571), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n570), .B1(KEYINPUT102), .B2(new_n571), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n604), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n609), .B2(new_n614), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n579), .A2(new_n584), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n577), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n573), .A2(KEYINPUT100), .A3(new_n574), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n639), .A2(new_n640), .B1(new_n580), .B2(new_n581), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n632), .B(new_n636), .C1(new_n641), .C2(new_n604), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  AND3_X1   g446(.A1(new_n635), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n643), .A2(KEYINPUT103), .A3(new_n634), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n643), .B2(new_n634), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n635), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n628), .A2(new_n654), .ZN(new_n655));
  NOR4_X1   g454(.A1(new_n492), .A2(new_n493), .A3(new_n559), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n439), .A2(new_n440), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n450), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n292), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n467), .A2(KEYINPUT40), .B1(new_n364), .B2(new_n366), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n464), .A2(new_n465), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n481), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n482), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n490), .A2(new_n489), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n485), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n559), .B1(new_n659), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n655), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT104), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n656), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n446), .A2(new_n373), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g475(.A(new_n660), .B1(new_n656), .B2(new_n671), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT105), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n679), .B(new_n660), .C1(new_n656), .C2(new_n671), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(G8gat), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n678), .B2(new_n680), .ZN(new_n685));
  OAI221_X1 g484(.A(new_n681), .B1(new_n677), .B2(new_n683), .C1(new_n685), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g485(.A(new_n487), .ZN(new_n687));
  AOI21_X1  g486(.A(G15gat), .B1(new_n672), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n491), .A2(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n491), .A2(KEYINPUT106), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT107), .Z(new_n694));
  AOI21_X1  g493(.A(new_n688), .B1(new_n672), .B2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n672), .A2(new_n481), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n669), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n595), .A2(new_n626), .ZN(new_n700));
  INV_X1    g499(.A(new_n654), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n673), .A2(G29gat), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n626), .B(KEYINPUT108), .Z(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n559), .A3(new_n701), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n659), .A2(new_n668), .ZN(new_n710));
  INV_X1    g509(.A(new_n595), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n710), .A2(new_n711), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g515(.A(new_n595), .B(new_n714), .C1(new_n659), .C2(new_n668), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n674), .B(new_n709), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n709), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n715), .A2(new_n713), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n492), .B2(new_n595), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(KEYINPUT110), .A3(new_n674), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n726), .A3(G29gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n707), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n707), .A2(new_n727), .A3(KEYINPUT111), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1328gat));
  INV_X1    g531(.A(G36gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n704), .A2(new_n733), .A3(new_n660), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n733), .B1(new_n725), .B2(new_n660), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n735), .A2(new_n736), .ZN(G1329gat));
  OAI211_X1 g536(.A(new_n692), .B(new_n709), .C1(new_n716), .C2(new_n717), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n487), .A2(G43gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n669), .A2(new_n702), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n669), .A2(KEYINPUT112), .A3(new_n702), .A4(new_n740), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT47), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  INV_X1    g547(.A(new_n491), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n709), .C1(new_n716), .C2(new_n717), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(G43gat), .B1(new_n743), .B2(new_n744), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n524), .B1(new_n725), .B2(new_n749), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n743), .A2(new_n744), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT47), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n747), .B1(new_n756), .B2(new_n746), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n753), .A2(new_n757), .ZN(G1330gat));
  AOI21_X1  g557(.A(new_n522), .B1(new_n725), .B2(new_n481), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n699), .A2(G50gat), .A3(new_n409), .A4(new_n703), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(KEYINPUT115), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n709), .B1(new_n716), .B2(new_n717), .ZN(new_n763));
  OAI21_X1  g562(.A(G50gat), .B1(new_n763), .B2(new_n409), .ZN(new_n764));
  INV_X1    g563(.A(new_n760), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n759), .A2(KEYINPUT114), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n761), .A2(new_n766), .B1(new_n767), .B2(KEYINPUT48), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT48), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT115), .B1(new_n759), .B2(new_n760), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n764), .A2(new_n762), .A3(new_n765), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n773), .ZN(G1331gat));
  NOR4_X1   g573(.A1(new_n492), .A2(new_n558), .A3(new_n627), .A4(new_n654), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n674), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT116), .B(G57gat), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1332gat));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n660), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT49), .B(G64gat), .Z(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(G1333gat));
  AOI21_X1  g581(.A(new_n599), .B1(new_n775), .B2(new_n692), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n487), .A2(G71gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n481), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n558), .A2(new_n626), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n710), .A2(new_n711), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n566), .A3(new_n674), .A4(new_n701), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n716), .A2(new_n717), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n701), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n673), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n566), .B2(new_n796), .ZN(G1336gat));
  NAND4_X1  g596(.A1(new_n792), .A2(new_n567), .A3(new_n660), .A4(new_n701), .ZN(new_n798));
  INV_X1    g597(.A(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n716), .B2(new_n717), .ZN(new_n800));
  OAI21_X1  g599(.A(G92gat), .B1(new_n800), .B2(new_n292), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n802), .B(new_n805), .ZN(G1337gat));
  INV_X1    g605(.A(G99gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n807), .A3(new_n687), .A4(new_n701), .ZN(new_n808));
  OAI21_X1  g607(.A(G99gat), .B1(new_n800), .B2(new_n691), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1338gat));
  OAI211_X1 g609(.A(new_n481), .B(new_n799), .C1(new_n716), .C2(new_n717), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT53), .B1(new_n812), .B2(KEYINPUT118), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n409), .A2(G106gat), .A3(new_n654), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n792), .A2(new_n814), .B1(new_n811), .B2(G106gat), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n813), .B(new_n815), .ZN(G1339gat));
  NOR2_X1   g615(.A1(new_n655), .A2(new_n558), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT103), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n644), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n649), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n643), .B2(new_n634), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n638), .A2(G230gat), .A3(new_n642), .A4(G233gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n647), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n498), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n544), .B2(new_n549), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n557), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n595), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT119), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n821), .A2(new_n824), .A3(new_n833), .A4(KEYINPUT55), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n648), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n829), .A2(new_n654), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n824), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n551), .A2(new_n557), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n595), .B1(new_n841), .B2(KEYINPUT120), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(new_n837), .C1(new_n835), .C2(new_n840), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n836), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n708), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n817), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n673), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n444), .A2(new_n436), .A3(new_n409), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(new_n292), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n558), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n487), .A2(new_n481), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n660), .A2(new_n673), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n847), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT121), .Z(new_n857));
  NOR2_X1   g656(.A1(new_n559), .A2(new_n311), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(G1340gat));
  AOI21_X1  g658(.A(G120gat), .B1(new_n850), .B2(new_n701), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n654), .A2(new_n313), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n857), .B2(new_n861), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n850), .A2(new_n863), .A3(new_n626), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n857), .A2(new_n708), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n863), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n660), .A2(new_n595), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n848), .A2(new_n867), .A3(new_n849), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT56), .Z(new_n870));
  AND2_X1   g669(.A1(new_n857), .A2(new_n711), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n867), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n749), .A2(new_n855), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT122), .B(new_n874), .C1(new_n847), .C2(new_n409), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n832), .A2(new_n834), .ZN(new_n876));
  INV_X1    g675(.A(new_n648), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n840), .ZN(new_n878));
  INV_X1    g677(.A(new_n837), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n595), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n626), .B1(new_n881), .B2(new_n836), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n481), .B1(new_n882), .B2(new_n817), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(new_n874), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n843), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n841), .A2(KEYINPUT120), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n595), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n708), .B1(new_n888), .B2(new_n836), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n481), .B1(new_n889), .B2(new_n817), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT122), .B1(new_n890), .B2(new_n874), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n873), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G141gat), .B1(new_n892), .B2(new_n559), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n692), .A2(new_n847), .A3(new_n409), .A4(new_n855), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n295), .A3(new_n558), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n893), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n883), .A2(KEYINPUT57), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n901), .A2(new_n701), .A3(new_n873), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G148gat), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n701), .B(new_n873), .C1(new_n885), .C2(new_n891), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n296), .A2(KEYINPUT59), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n296), .A3(new_n701), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n892), .B2(new_n846), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n300), .A3(new_n626), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n892), .B2(new_n595), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n692), .A2(new_n409), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(new_n301), .A3(new_n848), .A4(new_n868), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n674), .A2(new_n292), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n847), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(new_n849), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n558), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n847), .A2(new_n853), .A3(new_n923), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n559), .A2(new_n209), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n210), .A3(new_n701), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n927), .A2(new_n701), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n210), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT125), .Z(G1349gat));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n219), .A3(new_n626), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n927), .A2(new_n708), .ZN(new_n935));
  INV_X1    g734(.A(new_n224), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n925), .A2(new_n220), .A3(new_n711), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n927), .A2(new_n711), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G190gat), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n691), .A2(new_n922), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n890), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n558), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n945), .B(KEYINPUT126), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(new_n559), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n901), .A2(new_n902), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n947), .B1(new_n950), .B2(new_n952), .ZN(G1352gat));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n701), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n954), .B2(new_n948), .ZN(new_n955));
  NOR4_X1   g754(.A1(new_n945), .A2(new_n890), .A3(G204gat), .A4(new_n654), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n946), .A2(new_n261), .A3(new_n626), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n952), .A2(new_n626), .A3(new_n691), .A4(new_n922), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n946), .B2(new_n711), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n948), .A2(new_n260), .A3(new_n595), .ZN(new_n969));
  AOI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n969), .B2(new_n952), .ZN(G1355gat));
endmodule


