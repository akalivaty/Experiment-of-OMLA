

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  NAND2_X1 U325 ( .A1(n412), .A2(n411), .ZN(n414) );
  XNOR2_X1 U326 ( .A(n367), .B(n399), .ZN(n551) );
  INV_X1 U327 ( .A(KEYINPUT97), .ZN(n413) );
  XNOR2_X1 U328 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U329 ( .A(n414), .B(n413), .ZN(n460) );
  XNOR2_X1 U330 ( .A(n343), .B(n342), .ZN(n348) );
  XNOR2_X1 U331 ( .A(KEYINPUT26), .B(n403), .ZN(n568) );
  XOR2_X1 U332 ( .A(KEYINPUT38), .B(n452), .Z(n474) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U334 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XNOR2_X1 U335 ( .A(KEYINPUT100), .B(KEYINPUT36), .ZN(n310) );
  XOR2_X1 U336 ( .A(KEYINPUT75), .B(KEYINPUT64), .Z(n294) );
  XNOR2_X1 U337 ( .A(KEYINPUT11), .B(KEYINPUT76), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n309) );
  XOR2_X1 U339 ( .A(G99GAT), .B(G85GAT), .Z(n437) );
  XOR2_X1 U340 ( .A(G36GAT), .B(G190GAT), .Z(n371) );
  XOR2_X1 U341 ( .A(n437), .B(n371), .Z(n296) );
  XNOR2_X1 U342 ( .A(G218GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n302) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U345 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n434) );
  XOR2_X1 U347 ( .A(G134GAT), .B(n434), .Z(n300) );
  NAND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U351 ( .A(G50GAT), .B(G162GAT), .Z(n335) );
  XOR2_X1 U352 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n304) );
  XNOR2_X1 U353 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n335), .B(n305), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U357 ( .A(n309), .B(n308), .Z(n563) );
  INV_X1 U358 ( .A(n563), .ZN(n457) );
  XNOR2_X1 U359 ( .A(n310), .B(n457), .ZN(n583) );
  XOR2_X1 U360 ( .A(G78GAT), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U361 ( .A(G127GAT), .B(G71GAT), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U363 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n314) );
  XNOR2_X1 U364 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n325) );
  XNOR2_X1 U367 ( .A(G8GAT), .B(G183GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n317), .B(KEYINPUT77), .ZN(n370) );
  XOR2_X1 U369 ( .A(n370), .B(KEYINPUT78), .Z(n319) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U372 ( .A(KEYINPUT13), .B(G57GAT), .Z(n447) );
  XOR2_X1 U373 ( .A(n320), .B(n447), .Z(n323) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G1GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n321), .B(KEYINPUT70), .ZN(n433) );
  XOR2_X1 U376 ( .A(G22GAT), .B(G155GAT), .Z(n330) );
  XNOR2_X1 U377 ( .A(n433), .B(n330), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n579) );
  XOR2_X1 U380 ( .A(G204GAT), .B(KEYINPUT89), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT84), .B(KEYINPUT88), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n329) );
  INV_X1 U383 ( .A(KEYINPUT22), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n330), .B(KEYINPUT23), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U387 ( .A(n333), .B(KEYINPUT85), .Z(n343) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(G78GAT), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n334), .B(G148GAT), .ZN(n443) );
  XOR2_X1 U390 ( .A(n335), .B(n443), .Z(n337) );
  NAND2_X1 U391 ( .A1(G228GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U393 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n339) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n394) );
  XNOR2_X1 U396 ( .A(n394), .B(KEYINPUT24), .ZN(n340) );
  XOR2_X1 U397 ( .A(KEYINPUT86), .B(G218GAT), .Z(n345) );
  XNOR2_X1 U398 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U400 ( .A(G197GAT), .B(n346), .Z(n368) );
  INV_X1 U401 ( .A(n368), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n549) );
  XOR2_X1 U403 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U406 ( .A(G169GAT), .B(n351), .Z(n369) );
  XOR2_X1 U407 ( .A(KEYINPUT20), .B(G190GAT), .Z(n353) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G99GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U410 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n355) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n362) );
  XOR2_X1 U414 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XOR2_X1 U415 ( .A(G183GAT), .B(G176GAT), .Z(n359) );
  NAND2_X1 U416 ( .A1(G227GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n438), .B(n360), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n369), .B(n363), .ZN(n367) );
  XOR2_X1 U421 ( .A(KEYINPUT79), .B(G134GAT), .Z(n365) );
  XNOR2_X1 U422 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U424 ( .A(G113GAT), .B(n366), .ZN(n399) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n380) );
  XOR2_X1 U426 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U427 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n376) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G92GAT), .Z(n375) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n442) );
  XOR2_X1 U432 ( .A(n376), .B(n442), .Z(n378) );
  XNOR2_X1 U433 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n544) );
  INV_X1 U436 ( .A(n544), .ZN(n493) );
  NAND2_X1 U437 ( .A1(n551), .A2(n493), .ZN(n381) );
  NAND2_X1 U438 ( .A1(n549), .A2(n381), .ZN(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT25), .B(n382), .Z(n407) );
  XOR2_X1 U440 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n384) );
  XNOR2_X1 U441 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n398) );
  XOR2_X1 U443 ( .A(G155GAT), .B(G148GAT), .Z(n386) );
  XNOR2_X1 U444 ( .A(G29GAT), .B(G120GAT), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U446 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n388) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(G57GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U449 ( .A(n390), .B(n389), .Z(n396) );
  XOR2_X1 U450 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  NAND2_X1 U451 ( .A1(G225GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n547) );
  XOR2_X1 U457 ( .A(n544), .B(KEYINPUT27), .Z(n401) );
  XNOR2_X1 U458 ( .A(KEYINPUT94), .B(n401), .ZN(n502) );
  NOR2_X1 U459 ( .A1(n551), .A2(n549), .ZN(n402) );
  XOR2_X1 U460 ( .A(KEYINPUT95), .B(n402), .Z(n403) );
  NAND2_X1 U461 ( .A1(n502), .A2(n568), .ZN(n404) );
  XOR2_X1 U462 ( .A(KEYINPUT96), .B(n404), .Z(n405) );
  NOR2_X1 U463 ( .A1(n547), .A2(n405), .ZN(n406) );
  NAND2_X1 U464 ( .A1(n407), .A2(n406), .ZN(n412) );
  XNOR2_X1 U465 ( .A(KEYINPUT65), .B(KEYINPUT28), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n408), .B(n549), .ZN(n516) );
  NOR2_X1 U467 ( .A1(n551), .A2(n516), .ZN(n409) );
  NAND2_X1 U468 ( .A1(n502), .A2(n409), .ZN(n410) );
  NAND2_X1 U469 ( .A1(n410), .A2(n547), .ZN(n411) );
  NOR2_X1 U470 ( .A1(n579), .A2(n460), .ZN(n415) );
  NAND2_X1 U471 ( .A1(n583), .A2(n415), .ZN(n417) );
  INV_X1 U472 ( .A(KEYINPUT37), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n491) );
  XOR2_X1 U474 ( .A(G113GAT), .B(G36GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(G50GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U477 ( .A(G8GAT), .B(G197GAT), .Z(n421) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G22GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n428) );
  XOR2_X1 U481 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n425) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(KEYINPUT66), .B(n426), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U486 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n430) );
  XNOR2_X1 U487 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U489 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n570) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n451) );
  XOR2_X1 U493 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n440) );
  NAND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n441), .B(KEYINPUT73), .Z(n445) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U499 ( .A(n446), .B(KEYINPUT33), .Z(n449) );
  XNOR2_X1 U500 ( .A(n447), .B(KEYINPUT31), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n575) );
  OR2_X1 U503 ( .A1(n570), .A2(n575), .ZN(n462) );
  OR2_X1 U504 ( .A1(n491), .A2(n462), .ZN(n452) );
  NAND2_X1 U505 ( .A1(n474), .A2(n493), .ZN(n454) );
  XNOR2_X1 U506 ( .A(G36GAT), .B(KEYINPUT102), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(G1329GAT) );
  NAND2_X1 U508 ( .A1(n474), .A2(n551), .ZN(n456) );
  XNOR2_X1 U509 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n464) );
  INV_X1 U510 ( .A(n579), .ZN(n560) );
  NOR2_X1 U511 ( .A1(n457), .A2(n560), .ZN(n458) );
  XOR2_X1 U512 ( .A(KEYINPUT16), .B(n458), .Z(n459) );
  NOR2_X1 U513 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U514 ( .A(KEYINPUT98), .B(n461), .Z(n478) );
  NOR2_X1 U515 ( .A1(n478), .A2(n462), .ZN(n469) );
  NAND2_X1 U516 ( .A1(n469), .A2(n547), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(G1324GAT) );
  XOR2_X1 U518 ( .A(G8GAT), .B(KEYINPUT99), .Z(n466) );
  NAND2_X1 U519 ( .A1(n469), .A2(n493), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(G1325GAT) );
  XOR2_X1 U521 ( .A(G15GAT), .B(KEYINPUT35), .Z(n468) );
  NAND2_X1 U522 ( .A1(n469), .A2(n551), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(G1326GAT) );
  NAND2_X1 U524 ( .A1(n516), .A2(n469), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U526 ( .A1(n474), .A2(n547), .ZN(n473) );
  XNOR2_X1 U527 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT39), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(G1328GAT) );
  XOR2_X1 U530 ( .A(G50GAT), .B(KEYINPUT103), .Z(n476) );
  NAND2_X1 U531 ( .A1(n474), .A2(n516), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(G1331GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n480) );
  XNOR2_X1 U534 ( .A(n575), .B(KEYINPUT41), .ZN(n534) );
  XOR2_X1 U535 ( .A(KEYINPUT105), .B(n534), .Z(n554) );
  INV_X1 U536 ( .A(n554), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n570), .A2(n477), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n478), .A2(n490), .ZN(n485) );
  NAND2_X1 U539 ( .A1(n485), .A2(n547), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U541 ( .A(G57GAT), .B(n481), .Z(G1332GAT) );
  NAND2_X1 U542 ( .A1(n493), .A2(n485), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT106), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G64GAT), .B(n483), .ZN(G1333GAT) );
  NAND2_X1 U545 ( .A1(n551), .A2(n485), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n487) );
  NAND2_X1 U548 ( .A1(n485), .A2(n516), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n489) );
  XOR2_X1 U550 ( .A(G78GAT), .B(KEYINPUT108), .Z(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(G1335GAT) );
  NOR2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n497) );
  NAND2_X1 U553 ( .A1(n497), .A2(n547), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G85GAT), .B(n492), .ZN(G1336GAT) );
  XOR2_X1 U555 ( .A(G92GAT), .B(KEYINPUT109), .Z(n495) );
  NAND2_X1 U556 ( .A1(n497), .A2(n493), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1337GAT) );
  NAND2_X1 U558 ( .A1(n551), .A2(n497), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n501) );
  XOR2_X1 U561 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n499) );
  NAND2_X1 U562 ( .A1(n497), .A2(n516), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1339GAT) );
  NAND2_X1 U565 ( .A1(n547), .A2(n502), .ZN(n514) );
  NOR2_X1 U566 ( .A1(n570), .A2(n534), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(KEYINPUT46), .ZN(n504) );
  NOR2_X1 U568 ( .A1(n579), .A2(n504), .ZN(n505) );
  NAND2_X1 U569 ( .A1(n563), .A2(n505), .ZN(n506) );
  XNOR2_X1 U570 ( .A(KEYINPUT47), .B(n506), .ZN(n512) );
  XOR2_X1 U571 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n508) );
  NAND2_X1 U572 ( .A1(n579), .A2(n583), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U574 ( .A1(n509), .A2(n570), .ZN(n510) );
  NOR2_X1 U575 ( .A1(n575), .A2(n510), .ZN(n511) );
  NOR2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT48), .B(n513), .ZN(n543) );
  NOR2_X1 U578 ( .A1(n514), .A2(n543), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(KEYINPUT113), .ZN(n531) );
  NOR2_X1 U580 ( .A1(n516), .A2(n531), .ZN(n517) );
  NAND2_X1 U581 ( .A1(n517), .A2(n551), .ZN(n527) );
  NOR2_X1 U582 ( .A1(n570), .A2(n527), .ZN(n518) );
  XOR2_X1 U583 ( .A(KEYINPUT114), .B(n518), .Z(n519) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(n519), .ZN(G1340GAT) );
  NOR2_X1 U585 ( .A1(n527), .A2(n554), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n521) );
  XNOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1341GAT) );
  NOR2_X1 U590 ( .A1(n560), .A2(n527), .ZN(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(n526), .ZN(G1342GAT) );
  NOR2_X1 U594 ( .A1(n563), .A2(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(n530), .ZN(G1343GAT) );
  INV_X1 U598 ( .A(n531), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n532), .A2(n568), .ZN(n541) );
  NOR2_X1 U600 ( .A1(n570), .A2(n541), .ZN(n533) );
  XOR2_X1 U601 ( .A(G141GAT), .B(n533), .Z(G1344GAT) );
  NOR2_X1 U602 ( .A1(n541), .A2(n534), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n536) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1345GAT) );
  NOR2_X1 U607 ( .A1(n560), .A2(n541), .ZN(n539) );
  XOR2_X1 U608 ( .A(KEYINPUT120), .B(n539), .Z(n540) );
  XNOR2_X1 U609 ( .A(G155GAT), .B(n540), .ZN(G1346GAT) );
  NOR2_X1 U610 ( .A1(n563), .A2(n541), .ZN(n542) );
  XOR2_X1 U611 ( .A(G162GAT), .B(n542), .Z(G1347GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n567) );
  NAND2_X1 U616 ( .A1(n567), .A2(n549), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT55), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n562) );
  NOR2_X1 U619 ( .A1(n570), .A2(n562), .ZN(n553) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n553), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n562), .A2(n554), .ZN(n559) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n562), .ZN(n561) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n561), .Z(G1350GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G190GAT), .B(n566), .Z(G1351GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(n569), .Z(n574) );
  NOR2_X1 U635 ( .A1(n570), .A2(n574), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U640 ( .A(n574), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

