//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G137), .A3(new_n463), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n475), .B2(new_n461), .ZN(G160));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n463), .ZN(new_n477));
  OR3_X1    g052(.A1(new_n477), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(new_n477), .B2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n471), .A2(G2105), .A3(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n471), .A2(new_n461), .A3(new_n463), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n461), .A2(G102), .A3(G2104), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n471), .A2(G126), .A3(new_n463), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT68), .A2(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT68), .A2(G114), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(G2104), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n496), .A2(new_n502), .A3(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n461), .B1(new_n497), .B2(new_n500), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n518), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(G543), .A3(new_n517), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(G88), .B1(new_n526), .B2(G50), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n515), .A2(KEYINPUT71), .A3(G62), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(G62), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n514), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n527), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND2_X1  g111(.A1(new_n524), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n526), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n516), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n524), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n526), .A2(G52), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n514), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n526), .A2(G43), .B1(G651), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n524), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  INV_X1    g140(.A(G78), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n514), .A2(new_n565), .B1(new_n566), .B2(new_n510), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT73), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  OAI221_X1 g144(.A(new_n569), .B1(new_n566), .B2(new_n510), .C1(new_n514), .C2(new_n565), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G651), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n524), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n526), .A2(KEYINPUT9), .A3(G53), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n525), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n576), .ZN(G299));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NOR2_X1   g153(.A1(G168), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT74), .B1(new_n543), .B2(new_n544), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n579), .A2(new_n580), .ZN(G286));
  NAND2_X1  g156(.A1(new_n524), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n526), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT75), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n511), .A2(new_n513), .A3(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n522), .A2(G48), .A3(G543), .A4(new_n517), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n523), .ZN(G305));
  AOI22_X1  g167(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n516), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n524), .A2(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n526), .A2(G47), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n514), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n526), .A2(G54), .B1(G651), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT10), .B1(new_n523), .B2(new_n599), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g186(.A(KEYINPUT76), .B(G559), .Z(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(G860), .B2(new_n613), .ZN(G148));
  OAI21_X1  g189(.A(KEYINPUT77), .B1(new_n558), .B2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(KEYINPUT77), .B(new_n615), .S(new_n617), .Z(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n481), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n484), .A2(G123), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n622), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND4_X1  g200(.A1(new_n473), .A2(new_n461), .A3(new_n463), .A4(new_n465), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n625), .A2(new_n630), .ZN(G156));
  INV_X1    g206(.A(G14), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2438), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT81), .Z(new_n648));
  AOI211_X1 g223(.A(new_n632), .B(new_n648), .C1(new_n646), .C2(new_n643), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2100), .Z(new_n657));
  AND2_X1   g232(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  AOI21_X1  g234(.A(KEYINPUT18), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT82), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n662), .A2(new_n663), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT20), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n667), .A3(new_n670), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT22), .B(G1981), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G16), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT33), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1976), .ZN(new_n686));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT86), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT84), .B(G16), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT87), .B(G1971), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n686), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n699), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n481), .A2(G131), .ZN(new_n706));
  OR2_X1    g281(.A1(G95), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT83), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n484), .A2(G119), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G25), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n715), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n692), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(G290), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n692), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT85), .B(G1986), .Z(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NOR3_X1   g299(.A1(new_n718), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n705), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT36), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n705), .A2(new_n728), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n692), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n558), .B2(new_n692), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1341), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n735), .B2(KEYINPUT30), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(G28), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(KEYINPUT30), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G4), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n606), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1348), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n740), .B(new_n744), .C1(new_n713), .C2(new_n624), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n713), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n481), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n484), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n473), .A2(G105), .A3(new_n461), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  NAND4_X1  g326(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(new_n713), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G34), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(KEYINPUT24), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n713), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G160), .B2(new_n713), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n745), .B(new_n757), .C1(G2084), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G27), .A2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2078), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n713), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n713), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n713), .A2(G33), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n463), .A2(new_n465), .A3(G127), .ZN(new_n773));
  INV_X1    g348(.A(G115), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n464), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n481), .A2(KEYINPUT91), .A3(G139), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n779));
  INV_X1    g354(.A(G139), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n480), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n777), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT90), .B(KEYINPUT25), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n772), .B1(new_n787), .B2(new_n713), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G2072), .Z(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G21), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G168), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1966), .ZN(new_n792));
  MUX2_X1   g367(.A(G5), .B(G301), .S(G16), .Z(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT96), .Z(new_n794));
  AOI21_X1  g369(.A(new_n792), .B1(G1961), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n763), .A2(new_n771), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n794), .A2(G1961), .B1(G2084), .B2(new_n762), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n756), .B2(new_n755), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT97), .Z(new_n799));
  NAND2_X1  g374(.A1(G299), .A2(G16), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n692), .A2(KEYINPUT23), .A3(G20), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n802));
  INV_X1    g377(.A(G20), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n691), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n800), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT99), .B(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n796), .A2(new_n799), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n730), .A2(new_n731), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n713), .A2(G26), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n484), .A2(G128), .ZN(new_n811));
  OR2_X1    g386(.A1(G104), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n813));
  INV_X1    g388(.A(G140), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n811), .B(new_n813), .C1(new_n480), .C2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n810), .B1(new_n820), .B2(new_n713), .ZN(new_n821));
  MUX2_X1   g396(.A(new_n810), .B(new_n821), .S(KEYINPUT28), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2067), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n769), .A2(new_n770), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT98), .Z(new_n825));
  NOR3_X1   g400(.A1(new_n809), .A2(new_n823), .A3(new_n825), .ZN(G311));
  AND2_X1   g401(.A1(new_n730), .A2(new_n808), .ZN(new_n827));
  INV_X1    g402(.A(new_n823), .ZN(new_n828));
  INV_X1    g403(.A(new_n825), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n731), .ZN(G150));
  NAND2_X1  g405(.A1(new_n524), .A2(G93), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n526), .A2(G55), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n831), .B(new_n832), .C1(new_n516), .C2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT100), .Z(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT101), .B(G860), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n557), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n558), .A2(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT39), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n607), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n839), .B1(new_n846), .B2(new_n837), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT102), .Z(G145));
  INV_X1    g423(.A(G160), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n488), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n496), .A2(new_n502), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n820), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n819), .A2(new_n502), .A3(new_n496), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n752), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n752), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n787), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(new_n787), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n855), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n484), .A2(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  OAI221_X1 g440(.A(new_n862), .B1(new_n863), .B2(new_n864), .C1(new_n480), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n628), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n712), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n712), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n858), .A2(new_n861), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(KEYINPUT103), .A3(new_n870), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n858), .A2(new_n861), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n624), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n858), .A2(new_n861), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n624), .B1(new_n881), .B2(new_n873), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n851), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n877), .B1(new_n874), .B2(new_n876), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n873), .A3(new_n624), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n850), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g464(.A(new_n606), .B(G299), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n607), .A2(KEYINPUT104), .A3(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n890), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n894), .B2(KEYINPUT41), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT105), .B1(new_n890), .B2(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n842), .B(new_n616), .ZN(new_n900));
  MUX2_X1   g475(.A(new_n895), .B(new_n899), .S(new_n900), .Z(new_n901));
  XNOR2_X1  g476(.A(G303), .B(G288), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n721), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n901), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G868), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(G868), .B2(new_n835), .ZN(G295));
  OAI21_X1  g483(.A(new_n907), .B1(G868), .B2(new_n835), .ZN(G331));
  OAI21_X1  g484(.A(G171), .B1(new_n579), .B2(new_n580), .ZN(new_n910));
  NAND2_X1  g485(.A1(G168), .A2(G301), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n842), .ZN(new_n913));
  INV_X1    g488(.A(new_n842), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n910), .A3(new_n911), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n910), .A3(KEYINPUT106), .A4(new_n911), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n894), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n913), .A2(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n899), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n919), .A2(new_n922), .A3(new_n904), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(G37), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n904), .B1(new_n919), .B2(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT43), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n904), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n890), .A2(KEYINPUT41), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT107), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(KEYINPUT41), .B2(new_n894), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n917), .A2(new_n918), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n913), .A2(new_n915), .A3(new_n895), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NOR4_X1   g509(.A1(new_n923), .A2(new_n933), .A3(new_n934), .A4(G37), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n924), .B2(new_n925), .ZN(new_n937));
  INV_X1    g512(.A(new_n919), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n927), .A3(new_n921), .ZN(new_n939));
  INV_X1    g514(.A(new_n933), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n934), .A4(new_n887), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n936), .B1(new_n943), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g519(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n945));
  AOI21_X1  g520(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR4_X1   g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n468), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT108), .B(G1384), .Z(new_n951));
  AOI21_X1  g526(.A(KEYINPUT45), .B1(new_n852), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT46), .Z(new_n956));
  INV_X1    g531(.A(G2067), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n819), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n753), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(new_n953), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT124), .B(KEYINPUT47), .Z(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT125), .Z(new_n962));
  XNOR2_X1  g537(.A(new_n960), .B(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n752), .B(new_n954), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n711), .B(new_n716), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n953), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(G290), .A2(G1986), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n953), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT48), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n717), .A3(new_n712), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(G2067), .B2(new_n819), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n963), .B(new_n972), .C1(new_n953), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n852), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n977), .B(new_n978), .C1(new_n505), .C2(new_n506), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n503), .A2(new_n507), .A3(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT50), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n950), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1961), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G2078), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT45), .B(new_n951), .C1(new_n505), .C2(new_n506), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n950), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n852), .A2(new_n951), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n988), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT121), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(G40), .A4(G160), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n475), .A2(new_n461), .ZN(new_n999));
  INV_X1    g574(.A(new_n468), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(G40), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT121), .B1(new_n952), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n993), .A2(G2078), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .A4(new_n991), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n987), .A2(new_n994), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G171), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n986), .A2(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n978), .B1(new_n505), .B2(new_n506), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT113), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(new_n988), .A3(new_n980), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n950), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n983), .A2(new_n988), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1010), .A2(KEYINPUT115), .A3(new_n950), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1003), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1007), .A2(G301), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1006), .A2(new_n1018), .A3(KEYINPUT54), .ZN(new_n1019));
  XOR2_X1   g594(.A(G305), .B(G1981), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT49), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G305), .B(G1981), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1009), .A2(new_n980), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n950), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(new_n1024), .A3(new_n1026), .A4(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n683), .A2(G1976), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1026), .A2(G8), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1026), .A2(G8), .A3(new_n1028), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1027), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n1035), .B(KEYINPUT55), .Z(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1001), .A2(new_n947), .ZN(new_n1038));
  NAND3_X1  g613(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n991), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n989), .ZN(new_n1041));
  INV_X1    g616(.A(G1971), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n982), .A2(new_n770), .A3(new_n950), .A4(new_n984), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1034), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1036), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1009), .A2(KEYINPUT50), .A3(new_n980), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n503), .A2(new_n507), .A3(new_n976), .A4(new_n978), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(new_n950), .A3(KEYINPUT114), .A4(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1050), .A2(new_n770), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n950), .A3(new_n1049), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1051), .A2(new_n1054), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1047), .B1(new_n1055), .B2(new_n1037), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1019), .A2(new_n1046), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n985), .A2(G2084), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1059));
  INV_X1    g634(.A(G1966), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(G168), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1037), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1061), .B2(G168), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1037), .B1(new_n1061), .B2(G168), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1057), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1016), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT115), .B1(new_n1010), .B2(new_n950), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1003), .ZN(new_n1070));
  NOR4_X1   g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1014), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n987), .A2(new_n994), .ZN(new_n1072));
  OAI21_X1  g647(.A(G171), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1007), .A2(G301), .A3(new_n1004), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT122), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1078));
  AND4_X1   g653(.A1(G301), .A2(new_n987), .A3(new_n994), .A4(new_n1004), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT122), .B(new_n1076), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT120), .B(G1341), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT58), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1025), .B2(new_n950), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1038), .A2(new_n1039), .A3(new_n991), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n988), .B2(new_n983), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1087), .B2(new_n954), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n1088), .B2(new_n557), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1041), .A2(G1996), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(new_n558), .C1(new_n1091), .C2(new_n1085), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1026), .A2(G2067), .ZN(new_n1093));
  INV_X1    g668(.A(G1348), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n985), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1089), .A2(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n985), .A2(new_n1094), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1093), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n606), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n606), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT117), .B(G1956), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n1052), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT118), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1040), .A2(new_n989), .A3(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1105), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1103), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1097), .A2(new_n1102), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1087), .A2(new_n1109), .B1(new_n1052), .B2(new_n1104), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1108), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(KEYINPUT119), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1103), .B(new_n1111), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1101), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1114), .A2(new_n1119), .B1(new_n1120), .B2(new_n1111), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1067), .A2(new_n1082), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1027), .A2(new_n1029), .A3(new_n683), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(G1981), .B2(G305), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(G8), .A3(new_n1026), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1045), .A2(new_n1036), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1034), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1026), .A2(new_n1024), .A3(G8), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1026), .A2(G8), .A3(new_n1028), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1130), .A2(new_n1021), .B1(KEYINPUT52), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(new_n1031), .C1(new_n1045), .C2(new_n1036), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n1133), .B2(KEYINPUT116), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1061), .A2(new_n1037), .A3(G286), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1034), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1136), .B(new_n1137), .C1(new_n1036), .C2(new_n1045), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1134), .A2(new_n1127), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n1056), .A3(new_n1046), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1129), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1128), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1122), .A2(new_n1123), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1123), .B1(new_n1122), .B2(new_n1142), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1065), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1078), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1063), .A2(new_n1148), .A3(new_n1066), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(new_n1056), .A3(new_n1046), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1143), .A2(new_n1144), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n969), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT110), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G290), .A2(G1986), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(new_n953), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT111), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n968), .A2(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT112), .Z(new_n1161));
  OAI21_X1  g736(.A(new_n975), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT126), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1164), .B(new_n975), .C1(new_n1153), .C2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(G401), .A2(G227), .ZN(new_n1168));
  AND2_X1   g742(.A1(new_n888), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n939), .A2(new_n925), .A3(new_n887), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1170), .A2(KEYINPUT43), .ZN(new_n1171));
  AOI211_X1 g745(.A(new_n459), .B(G229), .C1(new_n1171), .C2(new_n941), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1172), .A3(KEYINPUT127), .ZN(new_n1173));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n1174));
  OAI211_X1 g748(.A(G319), .B(new_n680), .C1(new_n937), .C2(new_n942), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n888), .A2(new_n1168), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1177), .ZN(G308));
  NAND2_X1  g752(.A1(new_n1169), .A2(new_n1172), .ZN(G225));
endmodule


