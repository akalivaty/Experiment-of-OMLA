//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  AND2_X1   g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT9), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(KEYINPUT89), .ZN(new_n205));
  NOR2_X1   g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT90), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT91), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n203), .A2(new_n206), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT21), .ZN(new_n213));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G155gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT92), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n215), .B(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G183gat), .B(G211gat), .Z(new_n219));
  XOR2_X1   g018(.A(new_n218), .B(new_n219), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(KEYINPUT87), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(KEYINPUT87), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT88), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n222), .B2(new_n227), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n212), .A2(KEYINPUT21), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n218), .B(new_n219), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT95), .ZN(new_n241));
  XNOR2_X1  g040(.A(G43gat), .B(G50gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT15), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n247));
  AOI21_X1  g046(.A(G36gat), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G29gat), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n249), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n242), .A2(KEYINPUT15), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(KEYINPUT15), .A3(new_n242), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT7), .ZN(new_n260));
  INV_X1    g059(.A(G99gat), .ZN(new_n261));
  INV_X1    g060(.A(G106gat), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT8), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT93), .B(G85gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n260), .B(new_n263), .C1(G92gat), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G99gat), .B(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G232gat), .A2(G233gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n258), .A2(new_n267), .B1(KEYINPUT41), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n256), .A2(new_n257), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT86), .B1(new_n271), .B2(KEYINPUT17), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT17), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n267), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n258), .B2(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT94), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n281), .B(new_n278), .C1(new_n272), .C2(new_n275), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n270), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n241), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n269), .A2(KEYINPUT41), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n270), .ZN(new_n291));
  INV_X1    g090(.A(new_n275), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n273), .B1(new_n258), .B2(new_n274), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n279), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n276), .A2(KEYINPUT94), .A3(new_n279), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n284), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI211_X1 g098(.A(new_n284), .B(new_n291), .C1(new_n295), .C2(new_n296), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n285), .A2(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n284), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n241), .A4(new_n289), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n240), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n231), .B1(new_n271), .B2(KEYINPUT17), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n292), .B2(new_n293), .ZN(new_n308));
  NAND2_X1  g107(.A1(G229gat), .A2(G233gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n231), .A2(new_n258), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT18), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n231), .B(new_n258), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n309), .B(KEYINPUT13), .Z(new_n314));
  AOI22_X1  g113(.A1(new_n311), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G141gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(G197gat), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT11), .B(G169gat), .Z(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n319), .B(KEYINPUT12), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n308), .A2(KEYINPUT18), .A3(new_n309), .A4(new_n310), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n315), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n315), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G230gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n212), .A2(new_n267), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n277), .B1(new_n209), .B2(new_n211), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n212), .A2(KEYINPUT10), .A3(new_n267), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G176gat), .B(G204gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT96), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n338), .B(KEYINPUT97), .Z(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n333), .B2(new_n334), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n306), .A2(new_n325), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT31), .B(G50gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G22gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n288), .ZN(new_n354));
  XNOR2_X1  g153(.A(G141gat), .B(G148gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n352), .B(new_n354), .C1(new_n355), .C2(KEYINPUT2), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(G148gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G141gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G155gat), .B(G162gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n352), .A2(KEYINPUT2), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n351), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g165(.A(G211gat), .ZN(new_n367));
  INV_X1    g166(.A(G218gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G211gat), .A2(G218gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(G211gat), .A2(G218gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373));
  AND2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374));
  OAI221_X1 g173(.A(new_n371), .B1(KEYINPUT22), .B2(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  OAI22_X1  g174(.A1(new_n373), .A2(new_n374), .B1(new_n372), .B2(KEYINPUT22), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NOR2_X1   g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n372), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT75), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G228gat), .ZN(new_n387));
  INV_X1    g186(.A(G233gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n376), .A2(new_n370), .A3(new_n369), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n375), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n365), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n386), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n385), .A2(new_n375), .A3(new_n382), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n351), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n362), .B1(new_n363), .B2(new_n361), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n356), .A2(KEYINPUT76), .A3(new_n364), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n395), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n398), .A2(new_n405), .B1(new_n406), .B2(new_n366), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n350), .B(new_n394), .C1(new_n407), .C2(new_n390), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n395), .B2(new_n351), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n386), .B1(new_n411), .B2(new_n404), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n393), .A2(new_n390), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n412), .A2(new_n389), .B1(new_n413), .B2(new_n386), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n350), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n410), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n394), .B1(new_n407), .B2(new_n390), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT79), .B1(new_n414), .B2(new_n350), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n349), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n417), .B1(new_n410), .B2(new_n415), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n421), .A3(new_n416), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n348), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT0), .ZN(new_n430));
  XOR2_X1   g229(.A(G57gat), .B(G85gat), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n402), .A2(KEYINPUT3), .A3(new_n403), .ZN(new_n433));
  INV_X1    g232(.A(G120gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G113gat), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G120gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442));
  AND2_X1   g241(.A1(G127gat), .A2(G134gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(G127gat), .A2(G134gat), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT70), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n441), .A2(new_n442), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .A4(new_n439), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT68), .B(G134gat), .ZN(new_n452));
  INV_X1    g251(.A(G127gat), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n437), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n444), .B1(new_n455), .B2(new_n442), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n365), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n397), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n433), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT77), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT77), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n433), .A2(new_n458), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n446), .A2(new_n450), .B1(new_n456), .B2(new_n454), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n459), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(KEYINPUT4), .A3(new_n459), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n467), .B1(new_n404), .B2(new_n466), .ZN(new_n475));
  INV_X1    g274(.A(new_n472), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n465), .A2(new_n471), .A3(new_n474), .A4(new_n472), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n432), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT6), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n432), .A3(new_n479), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n485), .B2(KEYINPUT78), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G8gat), .B(G36gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G226gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(new_n388), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(G169gat), .A2(G176gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G169gat), .B2(G176gat), .ZN(new_n500));
  INV_X1    g299(.A(G169gat), .ZN(new_n501));
  INV_X1    g300(.A(G176gat), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n498), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G183gat), .ZN(new_n506));
  INV_X1    g305(.A(G190gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT24), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(G183gat), .A3(G190gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n511), .B1(G190gat), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n508), .A2(new_n510), .B1(new_n506), .B2(new_n507), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n504), .B1(new_n518), .B2(new_n503), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n507), .B1(new_n506), .B2(KEYINPUT27), .ZN(new_n520));
  AND2_X1   g319(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n523), .B2(KEYINPUT27), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT65), .B1(new_n524), .B2(KEYINPUT28), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n513), .A2(KEYINPUT27), .A3(new_n514), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT27), .ZN(new_n527));
  AOI21_X1  g326(.A(G190gat), .B1(new_n527), .B2(G183gat), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(G183gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n506), .A2(KEYINPUT27), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT28), .B(new_n507), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n525), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n501), .A2(new_n502), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n539), .A2(KEYINPUT26), .A3(new_n497), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n506), .A2(new_n507), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n497), .A2(KEYINPUT26), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI221_X4 g342(.A(new_n496), .B1(new_n517), .B2(new_n519), .C1(new_n538), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n517), .A2(new_n519), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n538), .A2(KEYINPUT67), .A3(new_n543), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT67), .B1(new_n538), .B2(new_n543), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n495), .A2(KEYINPUT29), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n395), .B(new_n544), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n495), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n538), .A2(new_n543), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n549), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n406), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n493), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n554), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n395), .ZN(new_n558));
  INV_X1    g357(.A(new_n544), .ZN(new_n559));
  INV_X1    g358(.A(new_n545), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT67), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n529), .A2(new_n530), .ZN(new_n562));
  AOI211_X1 g361(.A(KEYINPUT65), .B(KEYINPUT28), .C1(new_n526), .C2(new_n528), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n507), .A2(KEYINPUT28), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n532), .A2(new_n533), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT66), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n543), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n561), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n538), .A2(KEYINPUT67), .A3(new_n543), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n560), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n549), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n406), .B(new_n559), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n492), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n576), .A3(KEYINPUT30), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n558), .A2(new_n578), .A3(new_n492), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n428), .B1(new_n489), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n584));
  INV_X1    g383(.A(new_n475), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n472), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n469), .A2(new_n470), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n462), .B2(new_n464), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n588), .B2(new_n472), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n465), .A2(new_n471), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n584), .A3(new_n476), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n432), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n480), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT40), .A4(new_n432), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n593), .A2(new_n579), .A3(new_n577), .A4(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT80), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n596), .B1(new_n597), .B2(new_n406), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n559), .B1(new_n573), .B2(new_n574), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(KEYINPUT80), .A3(new_n395), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT81), .B1(new_n557), .B2(new_n395), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n551), .A2(new_n554), .A3(new_n603), .A4(new_n406), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT37), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n493), .A2(KEYINPUT37), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT38), .B1(new_n556), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n558), .A2(new_n575), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n493), .B1(new_n610), .B2(KEYINPUT37), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(new_n558), .B2(new_n575), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT38), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n481), .B(new_n576), .C1(new_n485), .C2(new_n480), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n427), .B(new_n595), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n548), .A2(new_n466), .ZN(new_n618));
  NAND2_X1  g417(.A1(G227gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n458), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT71), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT71), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n626), .A3(new_n623), .ZN(new_n627));
  XNOR2_X1  g426(.A(G15gat), .B(G43gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G71gat), .B(G99gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n622), .B2(KEYINPUT32), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n625), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n622), .B(KEYINPUT32), .C1(new_n623), .C2(new_n630), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n620), .B1(new_n618), .B2(new_n621), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT34), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT72), .ZN(new_n638));
  AOI211_X1 g437(.A(new_n620), .B(new_n638), .C1(new_n618), .C2(new_n621), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT73), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n636), .B2(new_n639), .ZN(new_n644));
  INV_X1    g443(.A(new_n638), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n646), .B(KEYINPUT73), .C1(new_n634), .C2(new_n635), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n632), .A2(new_n633), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT36), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n627), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n626), .B1(new_n622), .B2(new_n623), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n633), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n640), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT36), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n641), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n582), .A2(new_n617), .A3(new_n649), .A4(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT83), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT35), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n647), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n652), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n661), .A2(new_n427), .A3(new_n641), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n489), .A2(new_n581), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n481), .B1(new_n485), .B2(new_n480), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n427), .A2(new_n659), .A3(new_n580), .A4(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n640), .B1(new_n632), .B2(new_n633), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT82), .B1(new_n642), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT82), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n669), .A3(new_n641), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n657), .B(new_n658), .C1(new_n664), .C2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n580), .A3(new_n659), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n428), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n654), .A2(new_n669), .A3(new_n641), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n669), .B1(new_n654), .B2(new_n641), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n487), .B1(new_n483), .B2(new_n484), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n679), .A2(new_n680), .A3(new_n480), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n580), .B1(new_n681), .B2(new_n482), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n661), .A2(new_n427), .A3(new_n641), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT35), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n658), .B1(new_n685), .B2(new_n657), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n347), .B1(new_n673), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(KEYINPUT98), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(KEYINPUT98), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n489), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(new_n222), .ZN(G1324gat));
  INV_X1    g492(.A(new_n690), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n230), .B1(new_n694), .B2(new_n581), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G8gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n581), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n695), .B1(new_n699), .B2(KEYINPUT42), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(KEYINPUT100), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT100), .B1(new_n698), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(G1325gat));
  NAND2_X1  g503(.A1(new_n649), .A2(new_n656), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G15gat), .B1(new_n690), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n668), .A2(new_n670), .ZN(new_n708));
  INV_X1    g507(.A(G15gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n690), .B2(new_n710), .ZN(G1326gat));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n694), .A2(new_n712), .A3(new_n428), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT101), .B1(new_n690), .B2(new_n427), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n715), .B(new_n717), .ZN(G1327gat));
  OAI21_X1  g517(.A(new_n657), .B1(new_n664), .B2(new_n671), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT83), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n305), .B1(new_n720), .B2(new_n672), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n240), .A2(new_n325), .A3(new_n346), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(G29gat), .A3(new_n691), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT45), .Z(new_n725));
  AOI21_X1  g524(.A(new_n305), .B1(new_n685), .B2(new_n657), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n721), .B2(KEYINPUT44), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n722), .B(KEYINPUT102), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G29gat), .B1(new_n731), .B2(new_n691), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n725), .A2(new_n732), .ZN(G1328gat));
  OAI21_X1  g532(.A(G36gat), .B1(new_n731), .B2(new_n580), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n723), .A2(G36gat), .A3(new_n580), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n738), .A2(new_n721), .A3(new_n708), .A4(new_n722), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n730), .A2(new_n705), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n744));
  OAI211_X1 g543(.A(KEYINPUT47), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(G43gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n740), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(G1330gat));
  NAND3_X1  g549(.A1(new_n730), .A2(G50gat), .A3(new_n428), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n723), .A2(new_n427), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(G50gat), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g553(.A(new_n325), .ZN(new_n755));
  INV_X1    g554(.A(new_n346), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n306), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n719), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n489), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT105), .B(G57gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1332gat));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n581), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT49), .B(G64gat), .Z(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(G1333gat));
  XOR2_X1   g564(.A(new_n708), .B(KEYINPUT106), .Z(new_n766));
  AOI21_X1  g565(.A(G71gat), .B1(new_n758), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n705), .A2(G71gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g569(.A1(new_n758), .A2(new_n428), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n240), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n726), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n726), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT108), .Z(new_n779));
  NOR3_X1   g578(.A1(new_n756), .A2(new_n691), .A3(new_n264), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n305), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT44), .B(new_n782), .C1(new_n673), .C2(new_n686), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n755), .A2(new_n240), .A3(new_n756), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT107), .A4(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n489), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n264), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n781), .A2(new_n791), .ZN(G1336gat));
  NOR3_X1   g591(.A1(new_n756), .A2(G92gat), .A3(new_n580), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n728), .A2(KEYINPUT110), .A3(new_n581), .A4(new_n785), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n783), .A2(new_n784), .A3(new_n581), .A4(new_n785), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n800), .A3(G92gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(new_n801), .A3(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n581), .A3(new_n789), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n794), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n807), .B1(new_n810), .B2(KEYINPUT52), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n795), .B1(new_n808), .B2(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(KEYINPUT109), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n811), .B2(new_n814), .ZN(G1337gat));
  NAND3_X1  g614(.A1(new_n708), .A2(new_n261), .A3(new_n346), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT112), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n779), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n788), .A2(new_n705), .A3(new_n789), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n261), .B2(new_n819), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n728), .A2(new_n428), .A3(new_n785), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n262), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n262), .A2(new_n778), .A3(new_n428), .A4(new_n346), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n788), .A2(new_n428), .A3(new_n789), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n829), .B2(G106gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(G1339gat));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n333), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n331), .A2(new_n332), .A3(new_n327), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n338), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n333), .A2(new_n832), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n343), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n839), .B(new_n842), .C1(new_n323), .C2(new_n324), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n315), .A2(new_n321), .A3(new_n322), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n313), .A2(new_n314), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n319), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n346), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n305), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n237), .A2(new_n239), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n839), .A2(new_n842), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n847), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n301), .B(new_n304), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n240), .A2(new_n305), .A3(new_n325), .A4(new_n756), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT114), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(KEYINPUT114), .A3(new_n855), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n691), .A2(new_n581), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n708), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n427), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT115), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n859), .A2(new_n864), .A3(new_n427), .A4(new_n861), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n863), .A2(G113gat), .A3(new_n755), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n859), .A2(new_n489), .A3(new_n580), .A4(new_n662), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n436), .B1(new_n867), .B2(new_n325), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(G1340gat));
  NAND4_X1  g668(.A1(new_n863), .A2(G120gat), .A3(new_n346), .A4(new_n865), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n434), .B1(new_n867), .B2(new_n756), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1341gat));
  AND3_X1   g675(.A1(new_n863), .A2(new_n240), .A3(new_n865), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n240), .A2(new_n453), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n877), .A2(new_n453), .B1(new_n867), .B2(new_n878), .ZN(G1342gat));
  NAND2_X1  g678(.A1(new_n782), .A2(new_n452), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n782), .A3(new_n865), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G134gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1343gat));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n854), .A2(KEYINPUT114), .A3(new_n855), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n886), .B(new_n428), .C1(new_n887), .C2(new_n856), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n706), .A2(new_n860), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n854), .A2(new_n855), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n428), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT118), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n888), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n755), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n427), .A2(new_n581), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n706), .A2(new_n899), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n691), .B(new_n900), .C1(new_n857), .C2(new_n858), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n325), .A2(G141gat), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n898), .A2(G141gat), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n894), .B2(new_n325), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT58), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n903), .A2(new_n904), .B1(new_n908), .B2(new_n909), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n901), .A2(new_n359), .A3(new_n346), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n359), .A2(KEYINPUT59), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n346), .ZN(new_n914));
  XNOR2_X1  g713(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT57), .B(new_n428), .C1(new_n887), .C2(new_n856), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n892), .A2(new_n886), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n890), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n346), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n911), .B1(new_n914), .B2(new_n921), .ZN(G1345gat));
  NAND4_X1  g721(.A1(new_n895), .A2(G155gat), .A3(new_n240), .A4(new_n897), .ZN(new_n923));
  INV_X1    g722(.A(new_n901), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n353), .B1(new_n924), .B2(new_n850), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n923), .A2(KEYINPUT121), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT121), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n901), .B2(new_n782), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n305), .A2(new_n288), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n913), .B2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n489), .A2(new_n580), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n766), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n859), .A2(new_n427), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n501), .A3(new_n325), .ZN(new_n935));
  INV_X1    g734(.A(new_n932), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n683), .B(new_n936), .C1(new_n857), .C2(new_n858), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n755), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n935), .A2(new_n938), .ZN(G1348gat));
  NOR3_X1   g738(.A1(new_n934), .A2(new_n502), .A3(new_n756), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n937), .A2(new_n346), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n502), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(KEYINPUT122), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT122), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1349gat));
  OAI211_X1 g744(.A(new_n937), .B(new_n240), .C1(new_n535), .C2(new_n536), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n515), .B1(new_n934), .B2(new_n850), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n507), .A3(new_n782), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n934), .A2(new_n305), .ZN(new_n951));
  XNOR2_X1  g750(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(G190gat), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n951), .B2(G190gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1351gat));
  AOI21_X1  g755(.A(new_n427), .B1(new_n857), .B2(new_n858), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n705), .A2(new_n936), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n755), .ZN(new_n961));
  INV_X1    g760(.A(new_n958), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n916), .B2(new_n917), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n755), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  XNOR2_X1  g764(.A(KEYINPUT124), .B(G204gat), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n756), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT125), .B1(new_n959), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n957), .A2(new_n971), .A3(new_n958), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT126), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n970), .A2(new_n972), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n346), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n967), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n974), .A2(new_n975), .A3(new_n978), .A4(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n960), .A2(new_n367), .A3(new_n240), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n963), .A2(new_n240), .ZN(new_n984));
  AND4_X1   g783(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n367), .B1(KEYINPUT127), .B2(new_n986), .ZN(new_n987));
  AOI22_X1  g786(.A1(new_n984), .A2(new_n987), .B1(new_n983), .B2(KEYINPUT63), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n982), .B1(new_n985), .B2(new_n988), .ZN(G1354gat));
  NAND3_X1  g788(.A1(new_n960), .A2(new_n368), .A3(new_n782), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n963), .A2(new_n782), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n990), .B1(new_n991), .B2(new_n368), .ZN(G1355gat));
endmodule


