//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT69), .B(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n463), .A3(G137), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n463), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n479), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n486), .B(new_n488), .C1(new_n476), .C2(new_n477), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n466), .A2(new_n463), .A3(new_n492), .A4(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n464), .B2(new_n465), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n471), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G2104), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n491), .A2(new_n493), .B1(new_n499), .B2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n510), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT75), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n521), .B(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n523), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(KEYINPUT76), .B(new_n520), .C1(new_n524), .C2(new_n528), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n509), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n530), .B1(new_n535), .B2(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n522), .B(new_n523), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT76), .B1(new_n538), .B2(new_n520), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G168));
  AND2_X1   g115(.A1(new_n535), .A2(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n516), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n519), .A2(G90), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(new_n535), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n508), .A2(G56), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n516), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(G81), .B2(new_n519), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n531), .A2(G53), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n561), .A2(new_n562), .B1(G91), .B2(new_n519), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n516), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n562), .A2(new_n564), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n531), .A2(KEYINPUT79), .A3(G53), .A4(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n563), .A2(new_n566), .A3(new_n568), .A4(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  OR2_X1    g148(.A1(new_n514), .A2(new_n517), .ZN(G303));
  NAND2_X1  g149(.A1(new_n519), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n531), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n510), .A2(new_n579), .B1(new_n512), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n516), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n586), .A2(new_n516), .B1(new_n510), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n532), .A2(new_n534), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n535), .A2(G54), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n508), .A2(new_n509), .A3(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n516), .B1(new_n596), .B2(KEYINPUT80), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(KEYINPUT80), .B2(new_n596), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G284));
  OAI21_X1  g177(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G321));
  NAND2_X1  g178(.A1(G299), .A2(new_n600), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n600), .ZN(G280));
  INV_X1    g181(.A(G860), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n599), .B1(G559), .B2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g184(.A1(new_n554), .A2(new_n600), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n599), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n466), .A2(new_n472), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  AOI22_X1  g194(.A1(G123), .A2(new_n479), .B1(new_n480), .B2(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT83), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n629), .A2(new_n630), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT84), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT16), .Z(new_n641));
  AND2_X1   g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n641), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n628), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n639), .A2(new_n641), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n639), .A2(new_n641), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n627), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  OAI21_X1  g224(.A(G14), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(KEYINPUT85), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(KEYINPUT85), .A3(new_n649), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n617), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n623), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT87), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  OR3_X1    g252(.A1(new_n669), .A2(new_n675), .A3(new_n672), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(G33), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT25), .Z(new_n690));
  AOI22_X1  g265(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(new_n463), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n480), .A2(G139), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT93), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n688), .B1(new_n695), .B2(G29), .ZN(new_n696));
  INV_X1    g271(.A(G2072), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n480), .A2(G141), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT95), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n479), .A2(G129), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT26), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n704), .A2(new_n705), .B1(G105), .B2(new_n472), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n687), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n687), .B2(G32), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G2078), .ZN(new_n714));
  NOR2_X1   g289(.A1(G164), .A2(new_n687), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G27), .B2(new_n687), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n698), .B(new_n717), .C1(new_n714), .C2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(new_n599), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G4), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1348), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G11), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(G28), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n687), .B1(new_n725), .B2(G28), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n724), .B1(new_n726), .B2(new_n727), .C1(new_n622), .C2(new_n687), .ZN(new_n728));
  INV_X1    g303(.A(G2067), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n687), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NOR2_X1   g306(.A1(G104), .A2(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT92), .Z(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n734));
  AOI22_X1  g309(.A1(G128), .A2(new_n479), .B1(new_n480), .B2(G140), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n728), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n687), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G2084), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n738), .B(new_n744), .C1(new_n729), .C2(new_n737), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n723), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n747), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n721), .A2(new_n722), .B1(new_n749), .B2(G1961), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n718), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n747), .A2(KEYINPUT88), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n747), .A2(KEYINPUT88), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G19), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n555), .B2(new_n754), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT91), .ZN(new_n757));
  INV_X1    g332(.A(G1341), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n752), .A2(G20), .A3(new_n753), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT23), .ZN(new_n762));
  INV_X1    g337(.A(G299), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n747), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1956), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n751), .A2(new_n759), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n754), .A2(G22), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G166), .B2(new_n754), .ZN(new_n769));
  INV_X1    g344(.A(G1971), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G6), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n584), .B2(G16), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT32), .B(G1981), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G23), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT89), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G288), .B2(new_n747), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n771), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT90), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT34), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  AOI22_X1  g360(.A1(G119), .A2(new_n479), .B1(new_n480), .B2(G131), .ZN(new_n786));
  OAI221_X1 g361(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G25), .B(new_n788), .S(G29), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT35), .B(G1991), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n754), .A2(G24), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n588), .B1(new_n535), .B2(G47), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n754), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1986), .Z(new_n795));
  NAND4_X1  g370(.A1(new_n784), .A2(new_n785), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT36), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n687), .A2(G35), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G162), .B2(new_n687), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT29), .Z(new_n800));
  INV_X1    g375(.A(G2090), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n747), .A2(G21), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G168), .B2(new_n747), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G1966), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n805), .A2(G1966), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n802), .A2(new_n803), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n711), .A2(new_n712), .B1(G2084), .B2(new_n743), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n749), .A2(G1961), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT96), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n696), .A2(new_n697), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n767), .A2(new_n797), .A3(new_n808), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n719), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n820), .A2(new_n516), .B1(new_n510), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n535), .B2(G55), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n554), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n549), .A3(new_n553), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n819), .B(new_n827), .Z(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n829), .A2(new_n607), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n823), .A2(new_n607), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT97), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n834), .ZN(G145));
  XOR2_X1   g410(.A(new_n622), .B(G160), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n484), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n736), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n491), .A2(new_n493), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n500), .A2(new_n505), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n708), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n491), .B2(new_n493), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n840), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n709), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n846), .A2(new_n849), .A3(new_n695), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n694), .B1(new_n846), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n479), .A2(G130), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT99), .Z(new_n853));
  OR2_X1    g428(.A1(new_n463), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n854), .A2(new_n856), .B1(new_n480), .B2(G142), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n788), .B(new_n615), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n850), .A2(new_n851), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n694), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n848), .A2(new_n709), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n845), .A2(new_n708), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n846), .A2(new_n849), .A3(new_n695), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n838), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n861), .B1(new_n850), .B2(new_n851), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n860), .A3(new_n867), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n837), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g450(.A(KEYINPUT104), .B1(new_n823), .B2(G868), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n827), .B(KEYINPUT100), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n611), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n719), .A2(new_n763), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n599), .A2(G299), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n879), .A2(KEYINPUT41), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n880), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  NAND2_X1  g462(.A1(G290), .A2(KEYINPUT101), .ZN(new_n888));
  INV_X1    g463(.A(G288), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n793), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n888), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(G303), .A2(KEYINPUT102), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g471(.A1(G166), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n895), .A2(G305), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G305), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n891), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n793), .A2(new_n890), .ZN(new_n903));
  OAI21_X1  g478(.A(G288), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n894), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n900), .A2(new_n905), .A3(new_n906), .A4(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT42), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n887), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n600), .B1(new_n887), .B2(new_n911), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n876), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(G295));
  AOI21_X1  g492(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g494(.A1(G168), .A2(new_n827), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n825), .B(new_n826), .C1(new_n537), .C2(new_n539), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n920), .A2(G171), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G171), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n886), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G301), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n881), .A2(new_n882), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n920), .A2(G171), .A3(new_n921), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n924), .A2(new_n929), .A3(KEYINPUT105), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n910), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n908), .A2(new_n909), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n924), .A3(new_n929), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n870), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n919), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n870), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n924), .B2(new_n929), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(KEYINPUT43), .A3(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n938), .A2(KEYINPUT44), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n937), .A3(new_n919), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n934), .A2(new_n937), .A3(new_n945), .A4(new_n919), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n939), .B2(new_n940), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n948), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT45), .B1(new_n844), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G125), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n468), .B1(new_n478), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n463), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(G40), .A3(new_n473), .A4(new_n470), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n708), .B(G1996), .Z(new_n960));
  XNOR2_X1  g535(.A(new_n736), .B(new_n729), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n788), .B(new_n790), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT107), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(G290), .B(G1986), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n959), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G1384), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(G164), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n499), .A2(new_n506), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n841), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(KEYINPUT112), .A3(new_n971), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n970), .B1(new_n847), .B2(G1384), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n973), .A2(new_n976), .A3(new_n957), .A4(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n979));
  INV_X1    g554(.A(G1966), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n847), .A2(G1384), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n956), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n985));
  INV_X1    g560(.A(G2084), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n989));
  OAI21_X1  g564(.A(G8), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  NOR2_X1   g566(.A1(G168), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT51), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT123), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n990), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n978), .A2(new_n980), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n987), .A3(new_n981), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n992), .A2(KEYINPUT51), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT51), .B(G8), .C1(new_n1001), .C2(G286), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT122), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n996), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1001), .A2(new_n992), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n889), .A2(G1976), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n982), .A2(new_n957), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT110), .B1(new_n1015), .B2(G8), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1012), .B(new_n1014), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n584), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n581), .A2(new_n583), .A3(G1981), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1020), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1017), .A2(new_n1018), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1018), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1029), .A2(new_n1016), .B1(G1976), .B2(new_n889), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1019), .B(new_n1028), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n841), .B2(new_n974), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(KEYINPUT45), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT108), .B(new_n970), .C1(G164), .C2(G1384), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n956), .B1(new_n844), .B2(new_n971), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n770), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n984), .A2(new_n985), .A3(new_n801), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n1042));
  NAND3_X1  g617(.A1(G303), .A2(G8), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n1044));
  OAI22_X1  g619(.A1(G166), .A2(new_n991), .B1(KEYINPUT109), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1041), .A2(G8), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1032), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n975), .A2(new_n983), .A3(new_n950), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT50), .B1(new_n847), .B2(G1384), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n957), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1039), .B1(G2090), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1046), .B1(new_n1052), .B2(G8), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n984), .A2(new_n985), .ZN(new_n1056));
  INV_X1    g631(.A(G1961), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n951), .A2(new_n956), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2078), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n976), .A3(new_n973), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1035), .A2(new_n714), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT124), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1067), .A3(new_n1060), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1055), .A2(G301), .A3(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1010), .A2(new_n1011), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1073), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT115), .B(G1956), .Z(new_n1075));
  AND3_X1   g650(.A1(new_n1051), .A2(KEYINPUT116), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT116), .B1(new_n1051), .B2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n563), .A2(new_n568), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n566), .A2(new_n570), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1084));
  NOR2_X1   g659(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G299), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1078), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1056), .A2(new_n722), .ZN(new_n1092));
  NOR4_X1   g667(.A1(new_n956), .A2(new_n847), .A3(G1384), .A4(G2067), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT118), .B(new_n1093), .C1(new_n1056), .C2(new_n722), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n599), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1088), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(new_n1074), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1090), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1089), .A2(new_n1101), .A3(new_n1099), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1095), .A2(new_n1096), .B1(KEYINPUT60), .B2(new_n719), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n599), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT121), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT119), .B(G1996), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1015), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT58), .B(G1341), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1038), .A2(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1116), .B2(new_n555), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1116), .A2(new_n555), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g695(.A(new_n1108), .B1(KEYINPUT60), .B2(new_n719), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1110), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1100), .B1(new_n1104), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1061), .A2(G40), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n470), .A2(new_n473), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n463), .B1(new_n953), .B2(KEYINPUT125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n467), .A2(new_n1128), .A3(new_n468), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n847), .B2(new_n972), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1124), .B1(new_n1131), .B2(new_n951), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n844), .A2(new_n971), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n977), .A3(KEYINPUT126), .A4(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1961), .B1(new_n984), .B2(new_n985), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1064), .A2(new_n1067), .A3(new_n1060), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1067), .B1(new_n1064), .B2(new_n1060), .ZN(new_n1139));
  OAI211_X1 g714(.A(G301), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1069), .B2(G301), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1032), .A2(new_n1053), .A3(new_n1047), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1063), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1145), .B(G301), .C1(new_n1139), .C2(new_n1138), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1058), .A2(new_n1134), .A3(new_n1132), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1146), .B(KEYINPUT54), .C1(new_n1148), .C2(G301), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1143), .A2(new_n1144), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1072), .A2(new_n1123), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1047), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1024), .B(KEYINPUT111), .Z(new_n1153));
  NOR2_X1   g728(.A1(G288), .A2(G1976), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1028), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1152), .A2(new_n1032), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1001), .A2(G8), .A3(G168), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1055), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1041), .A2(G8), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT114), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1046), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1162), .B2(new_n1161), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1159), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(KEYINPUT63), .A4(new_n1048), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1157), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1151), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n968), .B1(new_n1071), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n958), .B1(new_n709), .B2(new_n961), .ZN(new_n1170));
  OR3_X1    g745(.A1(new_n958), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT46), .B1(new_n958), .B2(G1996), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT47), .Z(new_n1174));
  NOR2_X1   g749(.A1(G290), .A2(G1986), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n959), .A2(KEYINPUT48), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT48), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1175), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n958), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1176), .B(new_n1179), .C1(new_n965), .C2(new_n958), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n786), .A2(new_n790), .A3(new_n787), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n962), .A2(new_n1181), .B1(G2067), .B2(new_n736), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n959), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1174), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1169), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g760(.A1(G227), .A2(new_n461), .ZN(new_n1187));
  INV_X1    g761(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g762(.A(KEYINPUT127), .B1(G401), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  AND3_X1   g764(.A1(new_n648), .A2(KEYINPUT85), .A3(new_n649), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1191), .A2(new_n651), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1190), .B(new_n1187), .C1(new_n1192), .C2(new_n650), .ZN(new_n1193));
  NAND4_X1  g767(.A1(new_n1189), .A2(new_n874), .A3(new_n685), .A4(new_n1193), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n938), .A2(new_n941), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1195), .ZN(G308));
  INV_X1    g770(.A(G308), .ZN(G225));
endmodule


