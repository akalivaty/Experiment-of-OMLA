

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n560), .A2(n559), .ZN(G171) );
  OR2_X1 U554 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X2 U555 ( .A1(G2105), .A2(n532), .ZN(n884) );
  NOR2_X1 U556 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U557 ( .A1(G299), .A2(n693), .ZN(n694) );
  AND2_X1 U558 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U559 ( .A(n713), .B(KEYINPUT101), .ZN(n714) );
  INV_X1 U560 ( .A(KEYINPUT32), .ZN(n757) );
  NOR2_X1 U561 ( .A1(G651), .A2(n654), .ZN(n649) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U563 ( .A1(G91), .A2(n640), .ZN(n519) );
  XOR2_X1 U564 ( .A(KEYINPUT0), .B(G543), .Z(n654) );
  NAND2_X1 U565 ( .A1(G53), .A2(n649), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n523) );
  INV_X1 U567 ( .A(G651), .ZN(n524) );
  OR2_X1 U568 ( .A1(n524), .A2(n654), .ZN(n520) );
  XNOR2_X1 U569 ( .A(KEYINPUT65), .B(n520), .ZN(n643) );
  NAND2_X1 U570 ( .A1(n643), .A2(G78), .ZN(n521) );
  XOR2_X1 U571 ( .A(KEYINPUT70), .B(n521), .Z(n522) );
  NOR2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n528) );
  NOR2_X1 U573 ( .A1(G543), .A2(n524), .ZN(n526) );
  XNOR2_X1 U574 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n526), .B(n525), .ZN(n653) );
  NAND2_X1 U576 ( .A1(n653), .A2(G65), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(G299) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X2 U579 ( .A(KEYINPUT17), .B(n529), .Z(n885) );
  NAND2_X1 U580 ( .A1(n885), .A2(G138), .ZN(n536) );
  INV_X1 U581 ( .A(G2104), .ZN(n532) );
  AND2_X1 U582 ( .A1(n532), .A2(G2105), .ZN(n888) );
  NAND2_X1 U583 ( .A1(G126), .A2(n888), .ZN(n531) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U585 ( .A1(G114), .A2(n889), .ZN(n530) );
  AND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G102), .A2(n884), .ZN(n533) );
  AND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(G164) );
  NAND2_X1 U590 ( .A1(G101), .A2(n884), .ZN(n537) );
  XNOR2_X1 U591 ( .A(KEYINPUT23), .B(n537), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G125), .A2(n888), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G113), .A2(n889), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n885), .A2(G137), .ZN(n542) );
  AND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(G160) );
  XOR2_X1 U598 ( .A(G2443), .B(G2446), .Z(n545) );
  XNOR2_X1 U599 ( .A(G2427), .B(G2451), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n545), .B(n544), .ZN(n551) );
  XOR2_X1 U601 ( .A(G2430), .B(G2454), .Z(n547) );
  XNOR2_X1 U602 ( .A(G1348), .B(G1341), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U604 ( .A(G2435), .B(G2438), .Z(n548) );
  XNOR2_X1 U605 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U606 ( .A(n551), .B(n550), .Z(n552) );
  AND2_X1 U607 ( .A1(G14), .A2(n552), .ZN(G401) );
  NAND2_X1 U608 ( .A1(n649), .A2(G52), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n653), .A2(G64), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U611 ( .A1(n643), .A2(G77), .ZN(n555) );
  XOR2_X1 U612 ( .A(KEYINPUT69), .B(n555), .Z(n557) );
  NAND2_X1 U613 ( .A1(n640), .A2(G90), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G120), .ZN(G236) );
  INV_X1 U618 ( .A(G69), .ZN(G235) );
  INV_X1 U619 ( .A(G108), .ZN(G238) );
  INV_X1 U620 ( .A(G132), .ZN(G219) );
  INV_X1 U621 ( .A(G82), .ZN(G220) );
  NAND2_X1 U622 ( .A1(G88), .A2(n640), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G62), .A2(n653), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G75), .A2(n643), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G50), .A2(n649), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(G166) );
  NAND2_X1 U629 ( .A1(G63), .A2(n653), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G51), .A2(n649), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT6), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT75), .ZN(n577) );
  XNOR2_X1 U634 ( .A(KEYINPUT5), .B(KEYINPUT74), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n640), .A2(G89), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G76), .A2(n643), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n837) );
  NAND2_X1 U646 ( .A1(n837), .A2(G567), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT71), .ZN(n581) );
  XNOR2_X1 U648 ( .A(KEYINPUT11), .B(n581), .ZN(G234) );
  XOR2_X1 U649 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n583) );
  NAND2_X1 U650 ( .A1(G56), .A2(n653), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n583), .B(n582), .ZN(n590) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n640), .A2(G81), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G68), .A2(n643), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n588), .B(n587), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n649), .A2(G43), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n920) );
  INV_X1 U661 ( .A(G860), .ZN(n606) );
  OR2_X1 U662 ( .A1(n920), .A2(n606), .ZN(G153) );
  INV_X1 U663 ( .A(G171), .ZN(G301) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U665 ( .A1(G79), .A2(n643), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G54), .A2(n649), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G92), .A2(n640), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G66), .A2(n653), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT15), .ZN(n928) );
  INV_X1 U673 ( .A(G868), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n928), .A2(n602), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(G284) );
  NOR2_X1 U676 ( .A1(G286), .A2(n602), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT76), .ZN(n605) );
  NOR2_X1 U678 ( .A1(G299), .A2(G868), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n606), .A2(G559), .ZN(n607) );
  INV_X1 U681 ( .A(n928), .ZN(n906) );
  NAND2_X1 U682 ( .A1(n607), .A2(n906), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n920), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G868), .A2(n906), .ZN(n609) );
  NOR2_X1 U686 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G282) );
  XNOR2_X1 U688 ( .A(G2100), .B(KEYINPUT79), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G135), .A2(n885), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G111), .A2(n889), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G123), .A2(n888), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT18), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n615), .B(KEYINPUT77), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n884), .A2(G99), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n995) );
  XOR2_X1 U698 ( .A(G2096), .B(KEYINPUT78), .Z(n620) );
  XNOR2_X1 U699 ( .A(n995), .B(n620), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G559), .A2(n906), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(n920), .ZN(n664) );
  NOR2_X1 U703 ( .A1(G860), .A2(n664), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G67), .A2(n653), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G55), .A2(n649), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G80), .A2(n643), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G93), .A2(n640), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n667) );
  XNOR2_X1 U711 ( .A(n667), .B(KEYINPUT80), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n631), .B(n630), .ZN(G145) );
  NAND2_X1 U713 ( .A1(G60), .A2(n653), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G47), .A2(n649), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U716 ( .A(KEYINPUT68), .B(n634), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n643), .A2(G72), .ZN(n635) );
  XOR2_X1 U718 ( .A(KEYINPUT66), .B(n635), .Z(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(G85), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G86), .A2(n640), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G48), .A2(n649), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n653), .A2(G61), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G49), .A2(n649), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U734 ( .A1(G87), .A2(n654), .ZN(n655) );
  XOR2_X1 U735 ( .A(KEYINPUT81), .B(n655), .Z(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(G288) );
  XOR2_X1 U737 ( .A(G299), .B(G305), .Z(n658) );
  XNOR2_X1 U738 ( .A(G290), .B(n658), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n659) );
  XNOR2_X1 U740 ( .A(G288), .B(n659), .ZN(n660) );
  XOR2_X1 U741 ( .A(n661), .B(n660), .Z(n663) );
  XNOR2_X1 U742 ( .A(G166), .B(n667), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n909) );
  XNOR2_X1 U744 ( .A(n909), .B(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n665), .A2(G868), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n666), .B(KEYINPUT83), .ZN(n669) );
  NOR2_X1 U747 ( .A1(n667), .A2(G868), .ZN(n668) );
  NOR2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT84), .B(n670), .Z(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n675) );
  XNOR2_X1 U757 ( .A(KEYINPUT89), .B(n675), .ZN(n687) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U760 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G96), .A2(n678), .ZN(n841) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n841), .ZN(n679) );
  XNOR2_X1 U763 ( .A(KEYINPUT85), .B(n679), .ZN(n685) );
  NOR2_X1 U764 ( .A1(G235), .A2(G236), .ZN(n680) );
  XOR2_X1 U765 ( .A(KEYINPUT86), .B(n680), .Z(n681) );
  NOR2_X1 U766 ( .A1(G238), .A2(n681), .ZN(n682) );
  NAND2_X1 U767 ( .A1(G57), .A2(n682), .ZN(n842) );
  NAND2_X1 U768 ( .A1(G567), .A2(n842), .ZN(n683) );
  XNOR2_X1 U769 ( .A(KEYINPUT87), .B(n683), .ZN(n684) );
  NOR2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U771 ( .A(n686), .B(KEYINPUT88), .ZN(n844) );
  AND2_X1 U772 ( .A1(n687), .A2(n844), .ZN(n840) );
  NAND2_X1 U773 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  AND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n785) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n786) );
  NAND2_X1 U777 ( .A1(n785), .A2(n786), .ZN(n703) );
  XOR2_X1 U778 ( .A(KEYINPUT95), .B(n703), .Z(n719) );
  INV_X1 U779 ( .A(n719), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n696), .A2(G2072), .ZN(n689) );
  INV_X1 U781 ( .A(KEYINPUT27), .ZN(n688) );
  XNOR2_X1 U782 ( .A(n689), .B(n688), .ZN(n691) );
  XOR2_X1 U783 ( .A(G1956), .B(KEYINPUT97), .Z(n946) );
  NAND2_X1 U784 ( .A1(n946), .A2(n719), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U786 ( .A1(G299), .A2(n693), .ZN(n692) );
  XNOR2_X1 U787 ( .A(KEYINPUT28), .B(n692), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n694), .B(KEYINPUT100), .ZN(n701) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n703), .ZN(n695) );
  XNOR2_X1 U790 ( .A(KEYINPUT98), .B(n695), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n696), .A2(G2067), .ZN(n697) );
  XOR2_X1 U792 ( .A(KEYINPUT99), .B(n697), .Z(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n708) );
  NOR2_X1 U794 ( .A1(n928), .A2(n708), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n712) );
  INV_X1 U796 ( .A(n703), .ZN(n717) );
  INV_X1 U797 ( .A(n717), .ZN(n740) );
  INV_X1 U798 ( .A(G1996), .ZN(n972) );
  NOR2_X1 U799 ( .A1(n740), .A2(n972), .ZN(n702) );
  XOR2_X1 U800 ( .A(n702), .B(KEYINPUT26), .Z(n705) );
  NAND2_X1 U801 ( .A1(n703), .A2(G1341), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U803 ( .A1(n920), .A2(n706), .ZN(n707) );
  XNOR2_X1 U804 ( .A(n707), .B(KEYINPUT64), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n708), .A2(n928), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U808 ( .A(n716), .B(KEYINPUT29), .ZN(n750) );
  NOR2_X1 U809 ( .A1(n717), .A2(G1961), .ZN(n718) );
  XNOR2_X1 U810 ( .A(KEYINPUT94), .B(n718), .ZN(n722) );
  XOR2_X1 U811 ( .A(KEYINPUT25), .B(G2078), .Z(n976) );
  NOR2_X1 U812 ( .A1(n976), .A2(n719), .ZN(n720) );
  XNOR2_X1 U813 ( .A(KEYINPUT96), .B(n720), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n726) );
  NOR2_X1 U815 ( .A1(G301), .A2(n726), .ZN(n748) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n740), .ZN(n728) );
  AND2_X1 U817 ( .A1(G8), .A2(n728), .ZN(n723) );
  NAND2_X1 U818 ( .A1(G8), .A2(n740), .ZN(n784) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n784), .ZN(n729) );
  OR2_X1 U820 ( .A1(n723), .A2(n729), .ZN(n725) );
  OR2_X1 U821 ( .A1(n748), .A2(n725), .ZN(n724) );
  NOR2_X1 U822 ( .A1(n750), .A2(n724), .ZN(n738) );
  INV_X1 U823 ( .A(n725), .ZN(n736) );
  AND2_X1 U824 ( .A1(G301), .A2(n726), .ZN(n727) );
  XNOR2_X1 U825 ( .A(n727), .B(KEYINPUT102), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U827 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U828 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  NOR2_X1 U829 ( .A1(n732), .A2(G168), .ZN(n733) );
  NOR2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U831 ( .A(n735), .B(KEYINPUT31), .ZN(n752) );
  AND2_X1 U832 ( .A1(n736), .A2(n752), .ZN(n737) );
  NOR2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U834 ( .A(KEYINPUT103), .B(n739), .ZN(n760) );
  INV_X1 U835 ( .A(G8), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n784), .ZN(n742) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U838 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n743), .A2(G303), .ZN(n744) );
  NOR2_X1 U840 ( .A1(n745), .A2(n744), .ZN(n751) );
  AND2_X1 U841 ( .A1(G286), .A2(G8), .ZN(n746) );
  OR2_X1 U842 ( .A1(n751), .A2(n746), .ZN(n754) );
  INV_X1 U843 ( .A(n754), .ZN(n747) );
  OR2_X1 U844 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n756) );
  AND2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U848 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT104), .ZN(n762) );
  INV_X1 U851 ( .A(n762), .ZN(n773) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n926) );
  NOR2_X1 U854 ( .A1(n763), .A2(n926), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n773), .A2(n764), .ZN(n767) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n923) );
  INV_X1 U857 ( .A(n923), .ZN(n765) );
  NOR2_X1 U858 ( .A1(n784), .A2(n765), .ZN(n766) );
  AND2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U860 ( .A1(KEYINPUT33), .A2(n768), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n926), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U862 ( .A1(n769), .A2(n784), .ZN(n770) );
  NOR2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U864 ( .A(G1981), .B(G305), .Z(n933) );
  NAND2_X1 U865 ( .A1(n772), .A2(n933), .ZN(n780) );
  INV_X1 U866 ( .A(n773), .ZN(n776) );
  NAND2_X1 U867 ( .A1(G166), .A2(G8), .ZN(n774) );
  NOR2_X1 U868 ( .A1(G2090), .A2(n774), .ZN(n775) );
  XNOR2_X1 U869 ( .A(n777), .B(KEYINPUT105), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n778), .A2(n784), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n827) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XNOR2_X1 U873 ( .A(n781), .B(KEYINPUT24), .ZN(n782) );
  XNOR2_X1 U874 ( .A(n782), .B(KEYINPUT93), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n825) );
  INV_X1 U876 ( .A(n785), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT90), .B(n788), .Z(n829) );
  NAND2_X1 U879 ( .A1(G128), .A2(n888), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G116), .A2(n889), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U882 ( .A(n791), .B(KEYINPUT35), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G104), .A2(n884), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G140), .A2(n885), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U886 ( .A(KEYINPUT34), .B(n794), .Z(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U888 ( .A(n797), .B(KEYINPUT36), .ZN(n904) );
  XOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .Z(n798) );
  NOR2_X1 U890 ( .A1(n904), .A2(n798), .ZN(n1014) );
  NAND2_X1 U891 ( .A1(n904), .A2(n798), .ZN(n1001) );
  NOR2_X1 U892 ( .A1(n829), .A2(n1001), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT91), .B(n799), .Z(n831) );
  NAND2_X1 U894 ( .A1(G141), .A2(n885), .ZN(n801) );
  NAND2_X1 U895 ( .A1(G117), .A2(n889), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n884), .A2(G105), .ZN(n802) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n802), .Z(n803) );
  NOR2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n888), .A2(G129), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n882) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n882), .ZN(n1008) );
  NAND2_X1 U903 ( .A1(G1996), .A2(n882), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT92), .ZN(n815) );
  NAND2_X1 U905 ( .A1(G131), .A2(n885), .ZN(n809) );
  NAND2_X1 U906 ( .A1(G107), .A2(n889), .ZN(n808) );
  NAND2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U908 ( .A1(G95), .A2(n884), .ZN(n811) );
  NAND2_X1 U909 ( .A1(G119), .A2(n888), .ZN(n810) );
  NAND2_X1 U910 ( .A1(n811), .A2(n810), .ZN(n812) );
  OR2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n900) );
  NAND2_X1 U912 ( .A1(G1991), .A2(n900), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n1015) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n900), .ZN(n997) );
  NOR2_X1 U916 ( .A1(n816), .A2(n997), .ZN(n817) );
  NOR2_X1 U917 ( .A1(n1015), .A2(n817), .ZN(n818) );
  NOR2_X1 U918 ( .A1(n1008), .A2(n818), .ZN(n819) );
  XOR2_X1 U919 ( .A(KEYINPUT39), .B(n819), .Z(n820) );
  NOR2_X1 U920 ( .A1(n831), .A2(n820), .ZN(n821) );
  NOR2_X1 U921 ( .A1(n1014), .A2(n821), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n829), .A2(n822), .ZN(n823) );
  XOR2_X1 U923 ( .A(KEYINPUT106), .B(n823), .Z(n833) );
  INV_X1 U924 ( .A(n833), .ZN(n824) );
  OR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U926 ( .A1(n827), .A2(n826), .ZN(n835) );
  XNOR2_X1 U927 ( .A(G1986), .B(G290), .ZN(n930) );
  NOR2_X1 U928 ( .A1(n930), .A2(n1015), .ZN(n828) );
  NOR2_X1 U929 ( .A1(n829), .A2(n828), .ZN(n830) );
  OR2_X1 U930 ( .A1(n831), .A2(n830), .ZN(n832) );
  AND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U932 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U936 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n843), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U943 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U944 ( .A(KEYINPUT108), .B(n844), .ZN(G319) );
  XOR2_X1 U945 ( .A(G2096), .B(G2100), .Z(n846) );
  XNOR2_X1 U946 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U954 ( .A(G1981), .B(G1956), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1996), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U957 ( .A(G1986), .B(G1976), .Z(n856) );
  XNOR2_X1 U958 ( .A(G1961), .B(G1971), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U963 ( .A(G1991), .B(G2474), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U965 ( .A1(n888), .A2(G124), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G112), .A2(n889), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G100), .A2(n884), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G136), .A2(n885), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U973 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n870) );
  XNOR2_X1 U975 ( .A(n871), .B(n870), .ZN(n899) );
  NAND2_X1 U976 ( .A1(G130), .A2(n888), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G118), .A2(n889), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G106), .A2(n884), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G142), .A2(n885), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  XNOR2_X1 U983 ( .A(KEYINPUT110), .B(n877), .ZN(n878) );
  NOR2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U985 ( .A(G164), .B(n880), .Z(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n995), .B(n883), .ZN(n897) );
  NAND2_X1 U988 ( .A1(G103), .A2(n884), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G127), .A2(n888), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G115), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(KEYINPUT113), .B(n895), .Z(n1002) );
  XNOR2_X1 U997 ( .A(G160), .B(n1002), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n900), .B(G162), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(n904), .B(n903), .Z(n905) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n920), .B(KEYINPUT114), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(G171), .B(n906), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n909), .B(G286), .Z(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT116), .B(n917), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1020 ( .A(n920), .B(G1341), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(G299), .B(G1956), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(G1971), .B(KEYINPUT123), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n927), .B(G303), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(G1348), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(G1966), .B(G168), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT57), .B(n935), .Z(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G1961), .B(G171), .Z(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT122), .B(n940), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT56), .B(G16), .Z(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n1026) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n956) );
  XOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .Z(n945) );
  XNOR2_X1 U1042 ( .A(G4), .B(n945), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G20), .B(n946), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G1341), .B(G19), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G1981), .B(G6), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(KEYINPUT60), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n954), .B(KEYINPUT124), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1052 ( .A(KEYINPUT125), .B(n957), .Z(n965) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G1976), .B(G23), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1056 ( .A(KEYINPUT126), .B(n960), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G1986), .B(G24), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G5), .B(G1961), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1063 ( .A(KEYINPUT61), .B(n968), .Z(n969) );
  NOR2_X1 U1064 ( .A1(G16), .A2(n969), .ZN(n994) );
  INV_X1 U1065 ( .A(KEYINPUT55), .ZN(n1020) );
  XOR2_X1 U1066 ( .A(G34), .B(KEYINPUT121), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G2084), .B(KEYINPUT54), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(n971), .B(n970), .ZN(n985) );
  XNOR2_X1 U1069 ( .A(G32), .B(n972), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n973), .A2(G28), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(G2067), .B(G26), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(G33), .B(G2072), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n976), .B(G27), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(G1991), .B(G25), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n983), .B(KEYINPUT53), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1081 ( .A(G2090), .B(KEYINPUT120), .Z(n986) );
  XNOR2_X1 U1082 ( .A(G35), .B(n986), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(n1020), .B(n989), .ZN(n991) );
  INV_X1 U1085 ( .A(G29), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(G11), .A2(n992), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n1024) );
  XNOR2_X1 U1089 ( .A(G160), .B(G2084), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1092 ( .A(KEYINPUT117), .B(n999), .Z(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1013) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1002), .Z(n1004) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(KEYINPUT50), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1006), .B(KEYINPUT118), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1009), .Z(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT119), .B(n1018), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(G29), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1027), .Z(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

