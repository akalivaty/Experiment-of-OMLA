//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G238), .A3(G237), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT68), .Z(G261));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n453), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n479), .A2(KEYINPUT71), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n483), .A3(new_n462), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n463), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n489), .B1(new_n488), .B2(new_n487), .C1(G112), .C2(new_n462), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n464), .A2(new_n466), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(new_n462), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n464), .A3(new_n466), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n498), .A2(new_n464), .A3(new_n466), .A4(KEYINPUT74), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(KEYINPUT4), .A3(new_n502), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n468), .B2(new_n469), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(new_n462), .B2(G114), .ZN(new_n507));
  INV_X1    g082(.A(G102), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(new_n462), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n478), .A2(KEYINPUT73), .A3(G126), .A4(G2105), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n506), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OR3_X1    g096(.A1(new_n520), .A2(KEYINPUT75), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT75), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n517), .A2(new_n519), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G50), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NOR2_X1   g113(.A1(new_n528), .A2(new_n529), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n530), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n520), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n531), .A2(new_n547), .B1(new_n533), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G651), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n531), .A2(new_n554), .B1(new_n533), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n551), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n556), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  AOI22_X1  g146(.A1(new_n527), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n551), .ZN(new_n573));
  INV_X1    g148(.A(new_n531), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(G91), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n533), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n540), .A2(KEYINPUT9), .A3(G53), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(KEYINPUT78), .A3(new_n579), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n575), .A2(new_n582), .A3(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  NAND2_X1  g160(.A1(new_n574), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n540), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n527), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n551), .A2(new_n590), .B1(new_n591), .B2(new_n539), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n520), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n540), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n574), .A2(G85), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT80), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n540), .A2(G54), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n527), .A2(new_n530), .A3(G92), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  NOR2_X1   g190(.A1(new_n608), .A2(G559), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G860), .B2(new_n609), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(G148));
  NAND2_X1  g193(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n621));
  OAI21_X1  g196(.A(G868), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n491), .A2(KEYINPUT69), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n478), .A2(new_n467), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n473), .B(KEYINPUT70), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n492), .A2(G123), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT83), .Z(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n485), .A2(G135), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT85), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n645), .A2(new_n646), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n645), .A2(new_n646), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(G14), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT88), .ZN(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n664), .B(KEYINPUT17), .Z(new_n669));
  OAI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n662), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n665), .A3(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n685), .B1(KEYINPUT20), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(KEYINPUT20), .C2(new_n687), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1991), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1996), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n695), .B(new_n697), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  NOR2_X1   g274(.A1(G16), .A2(G21), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G168), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G28), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g278(.A(G29), .B1(new_n702), .B2(KEYINPUT30), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n701), .A2(G1966), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n485), .A2(G141), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  AOI22_X1  g283(.A1(G105), .A2(new_n628), .B1(new_n492), .B2(G129), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G29), .B2(G32), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n705), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G19), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n564), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1341), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n714), .B(new_n717), .C1(new_n712), .C2(new_n713), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT29), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G2090), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(G2090), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n725));
  INV_X1    g300(.A(G26), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(G29), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n482), .A2(G140), .A3(new_n484), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G116), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n463), .B1(new_n731), .B2(G2105), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n492), .A2(G128), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(new_n725), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G2067), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(G2067), .ZN(new_n738));
  NOR4_X1   g313(.A1(new_n723), .A2(new_n724), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G11), .ZN(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G4), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n609), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G1348), .ZN(new_n744));
  INV_X1    g319(.A(G2084), .ZN(new_n745));
  NAND2_X1  g320(.A1(G160), .A2(G29), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n746), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n744), .B1(new_n745), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G5), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G171), .B2(G16), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n638), .A2(G29), .B1(G1961), .B2(new_n757), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n758), .B1(G1961), .B2(new_n757), .C1(new_n743), .C2(G1348), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n701), .A2(G1966), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n755), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n718), .A2(new_n739), .A3(new_n740), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n719), .A2(G27), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G164), .B2(new_n719), .ZN(new_n764));
  MUX2_X1   g339(.A(new_n763), .B(new_n764), .S(KEYINPUT95), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2078), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n482), .A2(new_n484), .ZN(new_n769));
  INV_X1    g344(.A(G139), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n768), .B1(new_n769), .B2(new_n770), .C1(new_n771), .C2(new_n462), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n776));
  OAI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G33), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(G29), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2072), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n754), .A2(new_n745), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT94), .Z(new_n782));
  NOR4_X1   g357(.A1(new_n762), .A2(new_n766), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n719), .A2(G25), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n485), .A2(G131), .ZN(new_n785));
  OR2_X1    g360(.A1(G95), .A2(G2105), .ZN(new_n786));
  INV_X1    g361(.A(G107), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n463), .B1(new_n787), .B2(G2105), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n492), .A2(G119), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(new_n719), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n741), .A2(G24), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G290), .B2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n741), .A2(G22), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n741), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1971), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT32), .B(G1981), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT91), .B1(G16), .B2(G23), .ZN(new_n805));
  OR3_X1    g380(.A1(KEYINPUT91), .A2(G16), .A3(G23), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(G288), .C2(new_n741), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT33), .B(G1976), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n800), .A2(G1971), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n801), .A2(new_n804), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n798), .B1(KEYINPUT34), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n797), .A2(new_n795), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n812), .B(new_n813), .C1(KEYINPUT34), .C2(new_n811), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT36), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n741), .A2(G20), .ZN(new_n816));
  OAI211_X1 g391(.A(KEYINPUT23), .B(new_n816), .C1(new_n613), .C2(new_n741), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(KEYINPUT23), .B2(new_n816), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT96), .B(G1956), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n783), .A2(new_n815), .A3(new_n820), .ZN(G150));
  XNOR2_X1  g396(.A(G150), .B(KEYINPUT97), .ZN(G311));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n531), .A2(new_n823), .B1(new_n533), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n551), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n609), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n828), .B1(new_n561), .B2(new_n563), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n829), .A2(new_n562), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n831), .B1(new_n838), .B2(G860), .ZN(G145));
  XNOR2_X1  g414(.A(new_n495), .B(new_n790), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n729), .A2(new_n842), .A3(new_n733), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n729), .B2(new_n733), .ZN(new_n844));
  OAI21_X1  g419(.A(G164), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n734), .A2(KEYINPUT98), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n506), .A2(new_n514), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n729), .A2(new_n842), .A3(new_n733), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n710), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n845), .A2(new_n849), .A3(new_n710), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n841), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n773), .B1(new_n853), .B2(new_n774), .ZN(new_n854));
  INV_X1    g429(.A(new_n630), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n851), .B(new_n852), .C1(new_n841), .C2(new_n775), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n852), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT99), .B1(new_n858), .B2(new_n850), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n772), .B1(new_n859), .B2(KEYINPUT92), .ZN(new_n860));
  INV_X1    g435(.A(new_n856), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n630), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n638), .B(G160), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n492), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n864), .B1(new_n865), .B2(new_n866), .C1(new_n769), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n863), .B(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n857), .A2(new_n862), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n857), .B2(new_n862), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n840), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n869), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n860), .A2(new_n861), .A3(new_n630), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n840), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n857), .A2(new_n862), .A3(new_n869), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n872), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT100), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n872), .A2(new_n879), .A3(new_n883), .A4(new_n880), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT40), .B1(new_n882), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n609), .A2(new_n613), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n608), .A2(G299), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n837), .B1(new_n620), .B2(new_n621), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n608), .A2(G559), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT82), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(new_n619), .C1(new_n836), .C2(new_n835), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n891), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT101), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n608), .A2(G299), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n608), .A2(G299), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n892), .A3(new_n896), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(KEYINPUT101), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n898), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(G288), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n909));
  XOR2_X1   g484(.A(G303), .B(G305), .Z(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(KEYINPUT102), .A3(new_n910), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n907), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n920), .A2(new_n905), .A3(new_n898), .A4(new_n906), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G868), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n828), .A2(G868), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n888), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g501(.A(KEYINPUT103), .B(new_n924), .C1(new_n922), .C2(G868), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n925), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n913), .A2(new_n915), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n564), .A2(new_n829), .ZN(new_n932));
  INV_X1    g507(.A(new_n836), .ZN(new_n933));
  XNOR2_X1  g508(.A(G171), .B(G168), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(G171), .B(G286), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n835), .B2(new_n836), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n902), .A3(new_n903), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n935), .A2(new_n937), .A3(new_n890), .A4(new_n889), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(KEYINPUT104), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n931), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n913), .A2(new_n915), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT104), .B1(new_n939), .B2(new_n940), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n904), .B2(new_n938), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n949), .A3(new_n880), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n952), .B2(new_n931), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n946), .A2(new_n941), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n930), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n951), .C2(new_n956), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n950), .B2(KEYINPUT43), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n959), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n472), .A2(new_n964), .A3(new_n480), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n506), .B2(new_n514), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT111), .B(G8), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G288), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(G1976), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n971), .B(new_n972), .C1(G1976), .C2(new_n970), .ZN(new_n974));
  XNOR2_X1  g549(.A(G305), .B(G1981), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(G166), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(G303), .A2(G8), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n965), .B1(new_n966), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n847), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT112), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n966), .A2(new_n992), .A3(new_n987), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n847), .A2(new_n989), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n998), .A2(new_n965), .A3(new_n999), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n995), .A2(G2090), .B1(new_n1000), .B2(G1971), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n986), .B1(new_n1001), .B2(new_n968), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT62), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n965), .A3(new_n999), .ZN(new_n1004));
  INV_X1    g579(.A(G1966), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n479), .ZN(new_n1007));
  AOI22_X1  g582(.A1(G137), .A2(new_n1007), .B1(new_n628), .B2(G101), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n627), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1009));
  OAI211_X1 g584(.A(G40), .B(new_n1008), .C1(new_n1009), .C2(new_n462), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n990), .A2(KEYINPUT108), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n966), .A2(new_n1013), .A3(new_n987), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1011), .A2(new_n745), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G286), .A2(new_n968), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1006), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1006), .A2(new_n1015), .B1(G8), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1006), .A2(new_n1015), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(new_n968), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1003), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1000), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1028), .A3(KEYINPUT53), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1012), .A2(new_n1034), .A3(new_n965), .A4(new_n1014), .ZN(new_n1035));
  INV_X1    g610(.A(G1961), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G301), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1019), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(KEYINPUT51), .A3(new_n1017), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1024), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT62), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1025), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1023), .A2(new_n968), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G286), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1000), .A2(G1971), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1035), .A2(G2090), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n985), .A3(new_n984), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT63), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1045), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1002), .B1(new_n1043), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n980), .B1(new_n1055), .B2(new_n1053), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n978), .A2(new_n1057), .A3(new_n970), .ZN(new_n1058));
  OR2_X1    g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n969), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1045), .A3(new_n980), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1062), .B2(KEYINPUT63), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n994), .A2(G1956), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n1066));
  INV_X1    g641(.A(new_n580), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n575), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n998), .A2(new_n965), .A3(new_n999), .A4(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1064), .A2(new_n1065), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1069), .B(new_n1071), .C1(new_n994), .C2(G1956), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT113), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n967), .A2(G2067), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1035), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1078), .A2(new_n608), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1071), .B1(new_n994), .B2(G1956), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1069), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT114), .B(new_n1071), .C1(new_n994), .C2(G1956), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1075), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1087), .B(new_n1076), .C1(new_n1035), .C2(new_n1077), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT120), .B1(new_n1088), .B2(new_n608), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1090), .A3(new_n608), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1035), .A2(new_n1077), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1076), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n609), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n608), .A4(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT119), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1089), .A2(new_n1091), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1078), .A2(KEYINPUT60), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1085), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1105));
  INV_X1    g680(.A(new_n967), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT115), .B(KEYINPUT58), .Z(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(G1341), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1004), .A2(G1996), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n564), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1111), .B(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1105), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1072), .A2(new_n1074), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(KEYINPUT118), .A3(new_n1118), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1086), .B1(new_n1104), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1033), .A2(G301), .A3(new_n1037), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1126));
  AOI211_X1 g701(.A(KEYINPUT122), .B(new_n1030), .C1(new_n1000), .C2(new_n1026), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1037), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT54), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(new_n979), .ZN(new_n1131));
  NOR2_X1   g706(.A1(G301), .A2(KEYINPUT123), .ZN(new_n1132));
  OAI221_X1 g707(.A(KEYINPUT54), .B1(new_n1128), .B2(new_n1132), .C1(new_n1129), .C2(KEYINPUT123), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1002), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1053), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1056), .B(new_n1063), .C1(new_n1124), .C2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n998), .A2(new_n1010), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(G1996), .ZN(new_n1140));
  INV_X1    g715(.A(G2067), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n734), .B(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1138), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT106), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n790), .B(new_n793), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT107), .Z(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(G290), .B(G1986), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1138), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1137), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n791), .A2(new_n793), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1145), .A2(new_n1153), .B1(G2067), .B2(new_n734), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1138), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1138), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT46), .ZN(new_n1157));
  OR3_X1    g732(.A1(new_n1156), .A2(new_n1157), .A3(G1996), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1138), .B1(new_n1143), .B2(new_n1139), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1156), .B2(G1996), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT124), .B(KEYINPUT47), .Z(new_n1162));
  XNOR2_X1  g737(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1156), .A2(G1986), .A3(G290), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT48), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1155), .B(new_n1163), .C1(new_n1149), .C2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT125), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n1152), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g743(.A1(new_n660), .A2(G319), .A3(new_n678), .ZN(new_n1170));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g746(.A1(new_n660), .A2(new_n678), .A3(KEYINPUT126), .A4(G319), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n1175));
  AND3_X1   g749(.A1(new_n1174), .A2(new_n1175), .A3(new_n698), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1174), .B2(new_n698), .ZN(new_n1177));
  NOR2_X1   g751(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n954), .B1(new_n953), .B2(new_n949), .ZN(new_n1179));
  AND4_X1   g753(.A1(new_n954), .A2(new_n945), .A3(new_n880), .A4(new_n955), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g755(.A(new_n1178), .B(new_n1181), .C1(new_n882), .C2(new_n884), .ZN(G308));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n882), .B2(new_n884), .ZN(new_n1183));
  OAI21_X1  g757(.A(new_n1183), .B1(new_n1177), .B2(new_n1176), .ZN(G225));
endmodule


