

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(G2105), .A2(G2104), .ZN(n654) );
  NAND2_X1 U557 ( .A1(n762), .A2(G1341), .ZN(n725) );
  NOR2_X1 U558 ( .A1(n801), .A2(n800), .ZN(n543) );
  AND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  XNOR2_X1 U560 ( .A(n639), .B(KEYINPUT15), .ZN(n1002) );
  NOR2_X4 U561 ( .A1(n624), .A2(G2105), .ZN(n722) );
  OR2_X1 U562 ( .A1(n605), .A2(n604), .ZN(n1018) );
  AND2_X1 U563 ( .A1(n557), .A2(n529), .ZN(n554) );
  AND2_X1 U564 ( .A1(n538), .A2(n526), .ZN(n537) );
  NAND2_X1 U565 ( .A1(n536), .A2(n533), .ZN(n535) );
  NOR2_X1 U566 ( .A1(n1018), .A2(n726), .ZN(n727) );
  NOR2_X1 U567 ( .A1(n762), .A2(n979), .ZN(n724) );
  NAND2_X1 U568 ( .A1(G160), .A2(n723), .ZN(n762) );
  AND2_X1 U569 ( .A1(n819), .A2(G40), .ZN(n723) );
  OR2_X1 U570 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U571 ( .A1(n544), .A2(n527), .ZN(n548) );
  NOR2_X2 U572 ( .A1(n628), .A2(n627), .ZN(G160) );
  AND2_X1 U573 ( .A1(n546), .A2(n545), .ZN(n544) );
  XOR2_X2 U574 ( .A(KEYINPUT1), .B(n579), .Z(n612) );
  XNOR2_X2 U575 ( .A(KEYINPUT69), .B(n574), .ZN(n595) );
  NOR2_X1 U576 ( .A1(n559), .A2(n751), .ZN(n558) );
  NAND2_X1 U577 ( .A1(n556), .A2(n523), .ZN(n555) );
  NOR2_X1 U578 ( .A1(n767), .A2(n768), .ZN(n559) );
  INV_X1 U579 ( .A(n797), .ZN(n783) );
  NOR2_X1 U580 ( .A1(n783), .A2(KEYINPUT64), .ZN(n562) );
  INV_X1 U581 ( .A(G1384), .ZN(n547) );
  INV_X1 U582 ( .A(G286), .ZN(n556) );
  OR2_X1 U583 ( .A1(n774), .A2(n752), .ZN(n753) );
  NAND2_X1 U584 ( .A1(n554), .A2(n552), .ZN(n770) );
  NAND2_X1 U585 ( .A1(n553), .A2(n523), .ZN(n552) );
  XNOR2_X1 U586 ( .A(KEYINPUT94), .B(KEYINPUT32), .ZN(n769) );
  NAND2_X1 U587 ( .A1(n563), .A2(n561), .ZN(n560) );
  NOR2_X1 U588 ( .A1(n562), .A2(KEYINPUT33), .ZN(n561) );
  NOR2_X1 U589 ( .A1(n525), .A2(n566), .ZN(n546) );
  XNOR2_X1 U590 ( .A(n654), .B(n549), .ZN(n567) );
  INV_X1 U591 ( .A(KEYINPUT17), .ZN(n549) );
  NOR2_X1 U592 ( .A1(n833), .A2(n531), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n689) );
  XNOR2_X1 U594 ( .A(n551), .B(n550), .ZN(n626) );
  XNOR2_X1 U595 ( .A(KEYINPUT67), .B(KEYINPUT23), .ZN(n550) );
  NAND2_X1 U596 ( .A1(n722), .A2(G101), .ZN(n551) );
  AND2_X1 U597 ( .A1(n767), .A2(n768), .ZN(n523) );
  AND2_X1 U598 ( .A1(G286), .A2(KEYINPUT93), .ZN(n524) );
  AND2_X1 U599 ( .A1(G102), .A2(n722), .ZN(n525) );
  AND2_X1 U600 ( .A1(n737), .A2(n532), .ZN(n526) );
  NAND2_X1 U601 ( .A1(G126), .A2(n896), .ZN(n527) );
  XOR2_X1 U602 ( .A(n724), .B(KEYINPUT26), .Z(n528) );
  NAND2_X1 U603 ( .A1(n761), .A2(n760), .ZN(n772) );
  AND2_X1 U604 ( .A1(n558), .A2(n555), .ZN(n529) );
  INV_X1 U605 ( .A(KEYINPUT88), .ZN(n533) );
  AND2_X1 U606 ( .A1(n783), .A2(KEYINPUT64), .ZN(n530) );
  AND2_X1 U607 ( .A1(n1011), .A2(n845), .ZN(n531) );
  AND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n819) );
  INV_X1 U609 ( .A(KEYINPUT93), .ZN(n768) );
  NAND2_X1 U610 ( .A1(n534), .A2(n533), .ZN(n532) );
  INV_X1 U611 ( .A(n733), .ZN(n534) );
  NAND2_X1 U612 ( .A1(n537), .A2(n535), .ZN(n742) );
  INV_X1 U613 ( .A(n540), .ZN(n536) );
  NAND2_X1 U614 ( .A1(n540), .A2(n539), .ZN(n538) );
  AND2_X1 U615 ( .A1(n733), .A2(KEYINPUT88), .ZN(n539) );
  NAND2_X1 U616 ( .A1(n731), .A2(n730), .ZN(n540) );
  NAND2_X1 U617 ( .A1(n542), .A2(n541), .ZN(n848) );
  XNOR2_X1 U618 ( .A(n543), .B(KEYINPUT99), .ZN(n542) );
  NAND2_X1 U619 ( .A1(n567), .A2(G138), .ZN(n545) );
  INV_X1 U620 ( .A(n548), .ZN(G164) );
  INV_X1 U621 ( .A(n772), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n772), .A2(n524), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n564), .A2(n560), .ZN(n787) );
  NAND2_X1 U624 ( .A1(n565), .A2(n530), .ZN(n563) );
  NOR2_X1 U625 ( .A1(n565), .A2(KEYINPUT64), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n782), .B(KEYINPUT95), .ZN(n565) );
  AND2_X2 U627 ( .A1(n624), .A2(G2105), .ZN(n896) );
  AND2_X1 U628 ( .A1(G114), .A2(n897), .ZN(n566) );
  OR2_X1 U629 ( .A1(n785), .A2(n797), .ZN(n568) );
  INV_X1 U630 ( .A(G8), .ZN(n751) );
  OR2_X1 U631 ( .A1(n771), .A2(n751), .ZN(n752) );
  NOR2_X1 U632 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U633 ( .A1(n999), .A2(n568), .ZN(n786) );
  NAND2_X1 U634 ( .A1(n689), .A2(G89), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT4), .ZN(n576) );
  INV_X1 U636 ( .A(G651), .ZN(n578) );
  INV_X1 U637 ( .A(G543), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n570), .A2(KEYINPUT0), .ZN(n573) );
  INV_X1 U639 ( .A(KEYINPUT0), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n571), .A2(G543), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n580) );
  OR2_X1 U642 ( .A1(n578), .A2(n580), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G76), .A2(n595), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT5), .ZN(n585) );
  NOR2_X1 U646 ( .A1(G543), .A2(n578), .ZN(n579) );
  NAND2_X1 U647 ( .A1(G63), .A2(n612), .ZN(n582) );
  NOR2_X2 U648 ( .A1(G651), .A2(n580), .ZN(n684) );
  NAND2_X1 U649 ( .A1(G51), .A2(n684), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT6), .B(n583), .Z(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n586), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U654 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U655 ( .A1(G64), .A2(n612), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G52), .A2(n684), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G77), .A2(n595), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G90), .A2(n689), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U661 ( .A(KEYINPUT9), .B(n591), .Z(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(G171) );
  AND2_X1 U663 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U664 ( .A1(n689), .A2(G81), .ZN(n594) );
  XNOR2_X1 U665 ( .A(KEYINPUT12), .B(n594), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n595), .A2(G68), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(KEYINPUT72), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n600) );
  INV_X1 U669 ( .A(KEYINPUT13), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G56), .A2(n612), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n601), .Z(n603) );
  AND2_X1 U673 ( .A1(n684), .A2(G43), .ZN(n602) );
  INV_X1 U674 ( .A(G860), .ZN(n662) );
  OR2_X1 U675 ( .A1(n1018), .A2(n662), .ZN(G153) );
  INV_X1 U676 ( .A(G57), .ZN(G237) );
  INV_X1 U677 ( .A(G108), .ZN(G238) );
  NAND2_X1 U678 ( .A1(G75), .A2(n595), .ZN(n607) );
  NAND2_X1 U679 ( .A1(G88), .A2(n689), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U681 ( .A1(G62), .A2(n612), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G50), .A2(n684), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G166) );
  NAND2_X1 U685 ( .A1(G65), .A2(n612), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G53), .A2(n684), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT70), .B(n615), .Z(n619) );
  NAND2_X1 U689 ( .A1(G78), .A2(n595), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G91), .A2(n689), .ZN(n616) );
  AND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(G299) );
  INV_X1 U693 ( .A(G2104), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G125), .A2(n896), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n620), .B(KEYINPUT66), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G137), .A2(n567), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT68), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G113), .A2(n897), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G7), .A2(G661), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U703 ( .A(G567), .ZN(n717) );
  NOR2_X1 U704 ( .A1(G223), .A2(n717), .ZN(n630) );
  XOR2_X1 U705 ( .A(KEYINPUT71), .B(n630), .Z(n631) );
  XNOR2_X1 U706 ( .A(KEYINPUT11), .B(n631), .ZN(G234) );
  INV_X1 U707 ( .A(G171), .ZN(G301) );
  NAND2_X1 U708 ( .A1(G868), .A2(G301), .ZN(n641) );
  NAND2_X1 U709 ( .A1(G92), .A2(n689), .ZN(n638) );
  NAND2_X1 U710 ( .A1(G66), .A2(n612), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G79), .A2(n595), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G54), .A2(n684), .ZN(n634) );
  XNOR2_X1 U714 ( .A(KEYINPUT73), .B(n634), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  OR2_X1 U717 ( .A1(n1002), .A2(G868), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(G284) );
  INV_X1 U719 ( .A(G868), .ZN(n642) );
  NOR2_X1 U720 ( .A1(G286), .A2(n642), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n643), .B(KEYINPUT74), .ZN(n645) );
  NOR2_X1 U722 ( .A1(G299), .A2(G868), .ZN(n644) );
  NOR2_X1 U723 ( .A1(n645), .A2(n644), .ZN(G297) );
  NAND2_X1 U724 ( .A1(n662), .A2(G559), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n646), .A2(n1002), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n647), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U727 ( .A1(G868), .A2(n1018), .ZN(n650) );
  NAND2_X1 U728 ( .A1(G868), .A2(n1002), .ZN(n648) );
  NOR2_X1 U729 ( .A1(G559), .A2(n648), .ZN(n649) );
  NOR2_X1 U730 ( .A1(n650), .A2(n649), .ZN(G282) );
  NAND2_X1 U731 ( .A1(G123), .A2(n896), .ZN(n651) );
  XNOR2_X1 U732 ( .A(n651), .B(KEYINPUT18), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n722), .A2(G99), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n658) );
  XOR2_X1 U735 ( .A(KEYINPUT17), .B(n654), .Z(n893) );
  NAND2_X1 U736 ( .A1(G135), .A2(n893), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G111), .A2(n897), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n949) );
  XNOR2_X1 U740 ( .A(n949), .B(G2096), .ZN(n660) );
  INV_X1 U741 ( .A(G2100), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(G156) );
  NAND2_X1 U743 ( .A1(G559), .A2(n1002), .ZN(n661) );
  XOR2_X1 U744 ( .A(n1018), .B(n661), .Z(n698) );
  NAND2_X1 U745 ( .A1(n662), .A2(n698), .ZN(n669) );
  NAND2_X1 U746 ( .A1(G67), .A2(n612), .ZN(n664) );
  NAND2_X1 U747 ( .A1(G55), .A2(n684), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n664), .A2(n663), .ZN(n668) );
  NAND2_X1 U749 ( .A1(G80), .A2(n595), .ZN(n666) );
  NAND2_X1 U750 ( .A1(G93), .A2(n689), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n700) );
  XOR2_X1 U753 ( .A(n669), .B(n700), .Z(G145) );
  NAND2_X1 U754 ( .A1(G49), .A2(n684), .ZN(n671) );
  NAND2_X1 U755 ( .A1(G74), .A2(G651), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U757 ( .A1(n612), .A2(n672), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n580), .A2(G87), .ZN(n673) );
  NAND2_X1 U759 ( .A1(n674), .A2(n673), .ZN(G288) );
  NAND2_X1 U760 ( .A1(G73), .A2(n595), .ZN(n675) );
  XNOR2_X1 U761 ( .A(n675), .B(KEYINPUT2), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G61), .A2(n612), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G86), .A2(n689), .ZN(n676) );
  NAND2_X1 U764 ( .A1(n677), .A2(n676), .ZN(n680) );
  NAND2_X1 U765 ( .A1(G48), .A2(n684), .ZN(n678) );
  XNOR2_X1 U766 ( .A(KEYINPUT75), .B(n678), .ZN(n679) );
  NOR2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U768 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U769 ( .A(KEYINPUT76), .B(n683), .ZN(G305) );
  AND2_X1 U770 ( .A1(n595), .A2(G72), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G60), .A2(n612), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G47), .A2(n684), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n691) );
  NAND2_X1 U775 ( .A1(n689), .A2(G85), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n691), .A2(n690), .ZN(G290) );
  INV_X1 U777 ( .A(G299), .ZN(n738) );
  XNOR2_X1 U778 ( .A(KEYINPUT19), .B(KEYINPUT77), .ZN(n692) );
  XNOR2_X1 U779 ( .A(n692), .B(n700), .ZN(n693) );
  XNOR2_X1 U780 ( .A(n693), .B(G288), .ZN(n696) );
  XNOR2_X1 U781 ( .A(G166), .B(G305), .ZN(n694) );
  XNOR2_X1 U782 ( .A(n694), .B(G290), .ZN(n695) );
  XNOR2_X1 U783 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U784 ( .A(n738), .B(n697), .ZN(n921) );
  XNOR2_X1 U785 ( .A(n921), .B(n698), .ZN(n699) );
  NAND2_X1 U786 ( .A1(n699), .A2(G868), .ZN(n702) );
  OR2_X1 U787 ( .A1(G868), .A2(n700), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n702), .A2(n701), .ZN(G295) );
  NAND2_X1 U789 ( .A1(G2078), .A2(G2084), .ZN(n704) );
  XOR2_X1 U790 ( .A(KEYINPUT20), .B(KEYINPUT78), .Z(n703) );
  XNOR2_X1 U791 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n705), .A2(G2090), .ZN(n706) );
  XOR2_X1 U793 ( .A(KEYINPUT79), .B(n706), .Z(n707) );
  XNOR2_X1 U794 ( .A(KEYINPUT21), .B(n707), .ZN(n708) );
  NAND2_X1 U795 ( .A1(n708), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U796 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U797 ( .A1(G132), .A2(G82), .ZN(n709) );
  XNOR2_X1 U798 ( .A(n709), .B(KEYINPUT80), .ZN(n710) );
  XNOR2_X1 U799 ( .A(n710), .B(KEYINPUT22), .ZN(n711) );
  NOR2_X1 U800 ( .A1(G218), .A2(n711), .ZN(n712) );
  NAND2_X1 U801 ( .A1(G96), .A2(n712), .ZN(n854) );
  NAND2_X1 U802 ( .A1(G2106), .A2(n854), .ZN(n713) );
  XNOR2_X1 U803 ( .A(n713), .B(KEYINPUT81), .ZN(n719) );
  NAND2_X1 U804 ( .A1(G120), .A2(G69), .ZN(n714) );
  NOR2_X1 U805 ( .A1(G237), .A2(n714), .ZN(n715) );
  XOR2_X1 U806 ( .A(KEYINPUT82), .B(n715), .Z(n716) );
  NOR2_X1 U807 ( .A1(G238), .A2(n716), .ZN(n856) );
  NOR2_X1 U808 ( .A1(n717), .A2(n856), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(G319) );
  INV_X1 U810 ( .A(G319), .ZN(n721) );
  NAND2_X1 U811 ( .A1(G483), .A2(G661), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n853) );
  NAND2_X1 U813 ( .A1(n853), .A2(G36), .ZN(G176) );
  INV_X1 U814 ( .A(G166), .ZN(G303) );
  INV_X1 U815 ( .A(G1996), .ZN(n979) );
  NAND2_X1 U816 ( .A1(n528), .A2(n725), .ZN(n726) );
  XNOR2_X1 U817 ( .A(n727), .B(KEYINPUT65), .ZN(n731) );
  INV_X1 U818 ( .A(n762), .ZN(n746) );
  INV_X1 U819 ( .A(G1348), .ZN(n1026) );
  NOR2_X1 U820 ( .A1(n746), .A2(n1026), .ZN(n729) );
  INV_X1 U821 ( .A(G2067), .ZN(n974) );
  NOR2_X1 U822 ( .A1(n762), .A2(n974), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n1002), .A2(n732), .ZN(n730) );
  OR2_X1 U825 ( .A1(n1002), .A2(n732), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n746), .A2(G2072), .ZN(n734) );
  XNOR2_X1 U827 ( .A(n734), .B(KEYINPUT27), .ZN(n736) );
  INV_X1 U828 ( .A(G1956), .ZN(n1028) );
  NOR2_X1 U829 ( .A1(n1028), .A2(n746), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n737) );
  NOR2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U833 ( .A(n740), .B(KEYINPUT28), .Z(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U835 ( .A(KEYINPUT89), .B(KEYINPUT29), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n744), .B(n743), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n746), .A2(G1961), .ZN(n745) );
  XNOR2_X1 U838 ( .A(n745), .B(KEYINPUT87), .ZN(n748) );
  XNOR2_X1 U839 ( .A(KEYINPUT25), .B(G2078), .ZN(n973) );
  NAND2_X1 U840 ( .A1(n746), .A2(n973), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n755), .A2(G171), .ZN(n749) );
  NAND2_X1 U843 ( .A1(n750), .A2(n749), .ZN(n761) );
  NAND2_X1 U844 ( .A1(G8), .A2(n762), .ZN(n797) );
  NOR2_X1 U845 ( .A1(G1966), .A2(n797), .ZN(n774) );
  NOR2_X1 U846 ( .A1(G2084), .A2(n762), .ZN(n771) );
  XNOR2_X1 U847 ( .A(KEYINPUT30), .B(n753), .ZN(n754) );
  NOR2_X1 U848 ( .A1(G168), .A2(n754), .ZN(n758) );
  NOR2_X1 U849 ( .A1(G171), .A2(n755), .ZN(n756) );
  XNOR2_X1 U850 ( .A(n756), .B(KEYINPUT90), .ZN(n757) );
  XOR2_X1 U851 ( .A(KEYINPUT31), .B(n759), .Z(n760) );
  NOR2_X1 U852 ( .A1(G1971), .A2(n797), .ZN(n764) );
  NOR2_X1 U853 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U855 ( .A(n765), .B(KEYINPUT92), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n766), .A2(G303), .ZN(n767) );
  XNOR2_X1 U857 ( .A(n770), .B(n769), .ZN(n778) );
  NAND2_X1 U858 ( .A1(n771), .A2(G8), .ZN(n776) );
  XNOR2_X1 U859 ( .A(KEYINPUT91), .B(n772), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n788) );
  NOR2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  NOR2_X1 U864 ( .A1(G1971), .A2(G303), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n1006), .A2(n779), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n788), .A2(n780), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  NAND2_X1 U868 ( .A1(n781), .A2(n1007), .ZN(n782) );
  XOR2_X1 U869 ( .A(G1981), .B(G305), .Z(n784) );
  XNOR2_X1 U870 ( .A(KEYINPUT96), .B(n784), .ZN(n999) );
  NAND2_X1 U871 ( .A1(n1006), .A2(KEYINPUT33), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n801) );
  INV_X1 U873 ( .A(n788), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G8), .A2(G166), .ZN(n789) );
  NOR2_X1 U875 ( .A1(G2090), .A2(n789), .ZN(n790) );
  XOR2_X1 U876 ( .A(KEYINPUT97), .B(n790), .Z(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U878 ( .A(KEYINPUT98), .B(n793), .Z(n794) );
  NAND2_X1 U879 ( .A1(n794), .A2(n797), .ZN(n799) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U881 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  OR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G141), .A2(n893), .ZN(n803) );
  NAND2_X1 U885 ( .A1(G129), .A2(n896), .ZN(n802) );
  NAND2_X1 U886 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U887 ( .A1(n722), .A2(G105), .ZN(n804) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n804), .Z(n805) );
  NOR2_X1 U889 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U890 ( .A1(n897), .A2(G117), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n890) );
  NAND2_X1 U892 ( .A1(G1996), .A2(n890), .ZN(n809) );
  XNOR2_X1 U893 ( .A(n809), .B(KEYINPUT84), .ZN(n817) );
  NAND2_X1 U894 ( .A1(G131), .A2(n893), .ZN(n811) );
  NAND2_X1 U895 ( .A1(G119), .A2(n896), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U897 ( .A1(G95), .A2(n722), .ZN(n813) );
  NAND2_X1 U898 ( .A1(G107), .A2(n897), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U900 ( .A1(n815), .A2(n814), .ZN(n914) );
  NAND2_X1 U901 ( .A1(G1991), .A2(n914), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U903 ( .A(KEYINPUT85), .B(n818), .ZN(n960) );
  INV_X1 U904 ( .A(n960), .ZN(n821) );
  NAND2_X1 U905 ( .A1(G160), .A2(G40), .ZN(n820) );
  NOR2_X1 U906 ( .A1(n819), .A2(n820), .ZN(n845) );
  NAND2_X1 U907 ( .A1(n821), .A2(n845), .ZN(n834) );
  XNOR2_X1 U908 ( .A(G2067), .B(KEYINPUT37), .ZN(n842) );
  NAND2_X1 U909 ( .A1(G140), .A2(n893), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G104), .A2(n722), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U912 ( .A(KEYINPUT34), .B(n824), .ZN(n829) );
  NAND2_X1 U913 ( .A1(G128), .A2(n896), .ZN(n826) );
  NAND2_X1 U914 ( .A1(G116), .A2(n897), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U916 ( .A(n827), .B(KEYINPUT35), .Z(n828) );
  NOR2_X1 U917 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U918 ( .A(KEYINPUT36), .B(n830), .Z(n831) );
  XNOR2_X1 U919 ( .A(KEYINPUT83), .B(n831), .ZN(n904) );
  NOR2_X1 U920 ( .A1(n842), .A2(n904), .ZN(n958) );
  NAND2_X1 U921 ( .A1(n845), .A2(n958), .ZN(n840) );
  NAND2_X1 U922 ( .A1(n834), .A2(n840), .ZN(n832) );
  XNOR2_X1 U923 ( .A(n832), .B(KEYINPUT86), .ZN(n833) );
  XNOR2_X1 U924 ( .A(G1986), .B(G290), .ZN(n1011) );
  NOR2_X1 U925 ( .A1(G1996), .A2(n890), .ZN(n947) );
  INV_X1 U926 ( .A(n834), .ZN(n837) );
  NOR2_X1 U927 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U928 ( .A1(G1991), .A2(n914), .ZN(n950) );
  NOR2_X1 U929 ( .A1(n835), .A2(n950), .ZN(n836) );
  NOR2_X1 U930 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U931 ( .A1(n947), .A2(n838), .ZN(n839) );
  XNOR2_X1 U932 ( .A(KEYINPUT39), .B(n839), .ZN(n841) );
  NAND2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n844) );
  NAND2_X1 U934 ( .A1(n904), .A2(n842), .ZN(n843) );
  XNOR2_X1 U935 ( .A(n843), .B(KEYINPUT100), .ZN(n962) );
  NAND2_X1 U936 ( .A1(n844), .A2(n962), .ZN(n846) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U938 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U939 ( .A(n849), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U940 ( .A(G223), .ZN(n850) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U943 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U945 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U947 ( .A(G132), .ZN(G219) );
  INV_X1 U948 ( .A(G120), .ZN(G236) );
  INV_X1 U949 ( .A(G82), .ZN(G220) );
  INV_X1 U950 ( .A(G69), .ZN(G235) );
  INV_X1 U951 ( .A(n854), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n856), .A2(n855), .ZN(G261) );
  INV_X1 U953 ( .A(G261), .ZN(G325) );
  XOR2_X1 U954 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(G2072), .Z(n860) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U961 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1976), .B(G1961), .Z(n866) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1956), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(G1981), .B(G1966), .Z(n868) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U970 ( .A(KEYINPUT105), .B(G2474), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n874) );
  XOR2_X1 U972 ( .A(G1971), .B(KEYINPUT41), .Z(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G100), .A2(n722), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G112), .A2(n897), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(KEYINPUT106), .B(n877), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G124), .A2(n896), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n893), .A2(G136), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(G162) );
  NAND2_X1 U983 ( .A1(G130), .A2(n896), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G118), .A2(n897), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G142), .A2(n893), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G106), .A2(n722), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(G162), .B(n892), .ZN(n906) );
  NAND2_X1 U993 ( .A1(G139), .A2(n893), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G103), .A2(n722), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G127), .A2(n896), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n964) );
  XOR2_X1 U1001 ( .A(G160), .B(n964), .Z(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n917) );
  XOR2_X1 U1004 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT108), .B(KEYINPUT46), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n909), .B(KEYINPUT111), .Z(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT107), .B(KEYINPUT109), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n949), .B(n912), .Z(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1012 ( .A(G164), .B(n915), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G395) );
  XOR2_X1 U1015 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n920) );
  XNOR2_X1 U1016 ( .A(n1002), .B(G171), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n922), .B(n921), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n1018), .B(G286), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n925), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT114), .B(n926), .ZN(G397) );
  XOR2_X1 U1023 ( .A(KEYINPUT101), .B(KEYINPUT104), .Z(n928) );
  XNOR2_X1 U1024 ( .A(G1348), .B(G1341), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n928), .B(n927), .ZN(n938) );
  XOR2_X1 U1026 ( .A(G2427), .B(G2435), .Z(n930) );
  XNOR2_X1 U1027 ( .A(G2430), .B(G2438), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n930), .B(n929), .ZN(n934) );
  XOR2_X1 U1029 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n932) );
  XNOR2_X1 U1030 ( .A(G2446), .B(G2454), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(n932), .B(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(n934), .B(n933), .Z(n936) );
  XNOR2_X1 U1033 ( .A(G2451), .B(G2443), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n939), .A2(G14), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(G319), .A2(n945), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(G227), .A2(G229), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT49), .B(n940), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(G395), .A2(G397), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(G225) );
  INV_X1 U1043 ( .A(G225), .ZN(G308) );
  INV_X1 U1044 ( .A(G96), .ZN(G221) );
  INV_X1 U1045 ( .A(n945), .ZN(G401) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n948), .Z(n956) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1050 ( .A(KEYINPUT116), .B(n951), .Z(n954) );
  XNOR2_X1 U1051 ( .A(G2084), .B(G160), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT115), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT117), .B(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2072), .B(n964), .Z(n966) );
  XOR2_X1 U1060 ( .A(G164), .B(G2078), .Z(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1062 ( .A(KEYINPUT50), .B(n967), .Z(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT52), .B(n970), .ZN(n971) );
  INV_X1 U1065 ( .A(KEYINPUT55), .ZN(n995) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n995), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n972), .A2(G29), .ZN(n1059) );
  XNOR2_X1 U1068 ( .A(G2090), .B(G35), .ZN(n989) );
  XNOR2_X1 U1069 ( .A(n973), .B(G27), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n974), .B(G26), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G33), .B(G2072), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT118), .B(G32), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(n979), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT119), .B(n983), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(G28), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G25), .B(G1991), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(KEYINPUT120), .ZN(n993) );
  XOR2_X1 U1084 ( .A(G2084), .B(G34), .Z(n991) );
  XNOR2_X1 U1085 ( .A(KEYINPUT54), .B(n991), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(n995), .B(n994), .ZN(n997) );
  INV_X1 U1088 ( .A(G29), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(G11), .A2(n998), .ZN(n1057) );
  XNOR2_X1 U1091 ( .A(G16), .B(KEYINPUT56), .ZN(n1025) );
  XNOR2_X1 U1092 ( .A(G168), .B(G1966), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(n1001), .B(KEYINPUT57), .ZN(n1023) );
  XNOR2_X1 U1095 ( .A(n1002), .B(G1348), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(n1003), .B(KEYINPUT121), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(G1961), .B(G301), .ZN(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G166), .B(G1971), .ZN(n1013) );
  INV_X1 U1100 ( .A(n1006), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1102 ( .A(KEYINPUT122), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(G1956), .B(G299), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(G1341), .B(n1018), .Z(n1019) );
  XNOR2_X1 U1109 ( .A(KEYINPUT123), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1055) );
  INV_X1 U1113 ( .A(G16), .ZN(n1053) );
  XOR2_X1 U1114 ( .A(G1966), .B(G21), .Z(n1039) );
  XNOR2_X1 U1115 ( .A(KEYINPUT59), .B(G4), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(n1027), .B(n1026), .ZN(n1036) );
  XNOR2_X1 U1117 ( .A(G20), .B(n1028), .ZN(n1031) );
  XOR2_X1 U1118 ( .A(G1341), .B(G19), .Z(n1029) );
  XNOR2_X1 U1119 ( .A(KEYINPUT124), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(G6), .B(G1981), .ZN(n1032) );
  NOR2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1123 ( .A(n1034), .B(KEYINPUT125), .ZN(n1035) );
  NOR2_X1 U1124 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1125 ( .A(KEYINPUT60), .B(n1037), .ZN(n1038) );
  NAND2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1050) );
  XOR2_X1 U1127 ( .A(G1961), .B(G5), .Z(n1048) );
  XOR2_X1 U1128 ( .A(G1976), .B(G23), .Z(n1042) );
  XOR2_X1 U1129 ( .A(G22), .B(KEYINPUT126), .Z(n1040) );
  XNOR2_X1 U1130 ( .A(n1040), .B(G1971), .ZN(n1041) );
  NAND2_X1 U1131 ( .A1(n1042), .A2(n1041), .ZN(n1045) );
  XOR2_X1 U1132 ( .A(KEYINPUT127), .B(G1986), .Z(n1043) );
  XNOR2_X1 U1133 ( .A(G24), .B(n1043), .ZN(n1044) );
  NOR2_X1 U1134 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XNOR2_X1 U1135 ( .A(n1046), .B(KEYINPUT58), .ZN(n1047) );
  NAND2_X1 U1136 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NOR2_X1 U1137 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XNOR2_X1 U1138 ( .A(KEYINPUT61), .B(n1051), .ZN(n1052) );
  NAND2_X1 U1139 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  NAND2_X1 U1140 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  NOR2_X1 U1141 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NAND2_X1 U1142 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  XOR2_X1 U1143 ( .A(KEYINPUT62), .B(n1060), .Z(G311) );
  INV_X1 U1144 ( .A(G311), .ZN(G150) );
endmodule

