//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1326, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n205), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  AND2_X1   g0016(.A1(KEYINPUT64), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(KEYINPUT64), .A2(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n221), .A2(G50), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n205), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n216), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT75), .ZN(new_n247));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  AND2_X1   g0048(.A1(G1), .A2(G13), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n252), .B1(new_n251), .B2(new_n255), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n255), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(G226), .B2(new_n260), .ZN(new_n261));
  OR2_X1    g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1698), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G222), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(G1698), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n265), .B1(new_n266), .B2(new_n267), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n249), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT69), .B1(new_n249), .B2(new_n250), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G190), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n247), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n261), .A2(new_n275), .A3(KEYINPUT75), .A4(G190), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(new_n279), .B1(G200), .B2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n205), .B2(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n220), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT64), .ZN(new_n286));
  INV_X1    g0086(.A(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT64), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G33), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n288), .A2(KEYINPUT71), .A3(G33), .A4(new_n289), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g0094(.A(KEYINPUT8), .B(G58), .Z(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G150), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT72), .B1(new_n296), .B2(new_n298), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n285), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G1), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(G50), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n285), .B1(new_n304), .B2(G20), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n306), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n309), .B(KEYINPUT73), .Z(new_n310));
  NAND3_X1  g0110(.A1(new_n303), .A2(new_n310), .A3(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT9), .B1(new_n303), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT10), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n313), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n311), .A4(new_n280), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n276), .A2(G179), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n276), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n303), .A2(new_n310), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n295), .A2(new_n305), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n308), .B2(new_n295), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n288), .A2(new_n289), .ZN(new_n329));
  OAI211_X1 g0129(.A(KEYINPUT77), .B(new_n328), .C1(new_n329), .C2(new_n267), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT7), .A3(new_n287), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n219), .A2(new_n333), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT77), .B1(new_n336), .B2(new_n328), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n207), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n297), .A2(G159), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n285), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT7), .B1(new_n329), .B2(new_n267), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n333), .A2(new_n328), .A3(new_n287), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(G68), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n343), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n352), .B2(new_n344), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n327), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(G226), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n267), .A2(KEYINPUT78), .A3(G226), .A4(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  INV_X1    g0159(.A(G1698), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n267), .A2(G223), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n357), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n274), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n255), .A2(new_n364), .A3(G274), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT68), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(G232), .B2(new_n260), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(new_n277), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n260), .A2(G232), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n256), .B2(new_n257), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n274), .B2(new_n362), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(new_n372), .B2(G200), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n354), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n374), .B2(new_n376), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n320), .B1(new_n363), .B2(new_n368), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(G179), .B2(new_n372), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT18), .B1(new_n380), .B2(new_n354), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT79), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n328), .B1(new_n219), .B2(new_n333), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT7), .A4(G20), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n207), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n344), .B1(new_n385), .B2(new_n343), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n285), .ZN(new_n387));
  INV_X1    g0187(.A(new_n345), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n328), .B1(new_n329), .B2(new_n267), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n334), .A3(new_n330), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n326), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n363), .A2(new_n368), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G169), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n363), .A2(G179), .A3(new_n368), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n381), .A2(new_n382), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n382), .B1(new_n381), .B2(new_n400), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n378), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n366), .A2(new_n367), .B1(G238), .B2(new_n260), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G97), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(new_n360), .C1(new_n331), .C2(new_n332), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n274), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n405), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n405), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n415));
  INV_X1    g0215(.A(new_n273), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n271), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n408), .A2(new_n407), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n406), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n260), .A2(G238), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n256), .B2(new_n257), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT13), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n405), .A2(new_n410), .A3(new_n411), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(G179), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n423), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(G169), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n415), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT12), .B1(new_n305), .B2(G68), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n305), .A2(KEYINPUT12), .A3(G68), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n308), .A2(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n292), .A2(G77), .A3(new_n293), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT11), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n285), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n434), .B2(new_n285), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n428), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n422), .A2(G190), .A3(new_n423), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n425), .B2(G200), .ZN(new_n444));
  INV_X1    g0244(.A(G200), .ZN(new_n445));
  AOI211_X1 g0245(.A(KEYINPUT76), .B(new_n445), .C1(new_n422), .C2(new_n423), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n441), .B(new_n442), .C1(new_n444), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n258), .B1(G244), .B2(new_n260), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n267), .A2(G232), .A3(new_n360), .ZN(new_n449));
  INV_X1    g0249(.A(G107), .ZN(new_n450));
  OAI221_X1 g0250(.A(new_n449), .B1(new_n450), .B2(new_n267), .C1(new_n269), .C2(new_n208), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n274), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n320), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n294), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n295), .A2(new_n297), .B1(new_n329), .B2(G77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n285), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n305), .A2(G77), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n308), .B2(G77), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n454), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G179), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n448), .A2(new_n465), .A3(new_n452), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n453), .A2(G200), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n460), .A2(KEYINPUT74), .A3(new_n462), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT74), .B1(new_n460), .B2(new_n462), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n468), .B1(new_n277), .B2(new_n453), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n440), .A2(new_n447), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n324), .A2(new_n404), .A3(new_n472), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT85), .B(KEYINPUT22), .Z(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G87), .A3(new_n219), .A4(new_n267), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n219), .A2(new_n267), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n477), .B2(new_n209), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT23), .A2(G107), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(G20), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT23), .A2(G107), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n329), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n347), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT24), .A4(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n305), .B1(G1), .B2(new_n282), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n285), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n305), .A2(G107), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT25), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT86), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n210), .A2(G1698), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n331), .B2(new_n332), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n267), .A2(KEYINPUT87), .A3(new_n500), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G294), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n274), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n304), .A2(G45), .ZN(new_n509));
  OR2_X1    g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n251), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n259), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G264), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT88), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n507), .A2(new_n274), .B1(G264), .B2(new_n514), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT88), .B1(new_n519), .B2(new_n513), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n277), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n445), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n499), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n487), .A2(new_n486), .B1(new_n496), .B2(new_n497), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(new_n517), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n513), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(G169), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n516), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G179), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n524), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  AND2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n450), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n219), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n297), .A2(G77), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT81), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n450), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n532), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n541), .B(new_n538), .C1(new_n544), .C2(new_n219), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n348), .A2(G107), .A3(new_n349), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n540), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n285), .ZN(new_n548));
  OAI21_X1  g0348(.A(G97), .B1(new_n285), .B2(new_n489), .ZN(new_n549));
  INV_X1    g0349(.A(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n305), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  OAI211_X1 g0358(.A(G250), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(new_n360), .C1(new_n331), .C2(new_n332), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT4), .B1(new_n264), .B2(G244), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n274), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n254), .A2(G1), .ZN(new_n565));
  INV_X1    g0365(.A(new_n511), .ZN(new_n566));
  NOR2_X1   g0366(.A1(KEYINPUT5), .A2(G41), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G257), .A3(new_n364), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n513), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n320), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n513), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n513), .A3(KEYINPUT83), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n564), .A2(new_n574), .A3(new_n465), .A4(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n557), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n285), .A2(new_n547), .B1(new_n553), .B2(new_n555), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n564), .A2(new_n574), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n560), .A2(new_n561), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n558), .A4(new_n559), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n572), .B1(new_n583), .B2(new_n274), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G190), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n578), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n364), .A2(G274), .A3(new_n565), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n364), .A2(G250), .A3(new_n509), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G238), .B(new_n360), .C1(new_n331), .C2(new_n332), .ZN(new_n590));
  OAI211_X1 g0390(.A(G244), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G116), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI211_X1 g0393(.A(G179), .B(new_n589), .C1(new_n274), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n274), .A2(new_n593), .ZN(new_n595));
  INV_X1    g0395(.A(new_n589), .ZN(new_n596));
  AOI21_X1  g0396(.A(G169), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G13), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(G1), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n455), .A2(G20), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n490), .A2(new_n456), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n219), .A2(new_n267), .A3(G68), .ZN(new_n603));
  NAND3_X1  g0403(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n288), .A2(new_n289), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n534), .A2(new_n209), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n292), .A2(G97), .A3(new_n293), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n601), .B(new_n602), .C1(new_n611), .C2(new_n347), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n598), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n595), .A2(new_n277), .A3(new_n596), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n589), .B1(new_n274), .B2(new_n593), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(G200), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n609), .A2(new_n610), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n285), .B1(new_n617), .B2(new_n608), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n490), .A2(G87), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n601), .A4(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n577), .A2(new_n586), .A3(new_n613), .A4(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n600), .A2(G20), .B1(new_n304), .B2(G33), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n284), .A2(new_n220), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(G116), .A4(new_n283), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G116), .B2(new_n305), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n282), .A2(G97), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n219), .A2(new_n558), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G116), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G20), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n285), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n626), .A2(new_n558), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n219), .B1(G20), .B2(new_n628), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n285), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n625), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n514), .A2(G270), .B1(new_n251), .B2(new_n512), .ZN(new_n637));
  OAI211_X1 g0437(.A(G264), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n638));
  OAI211_X1 g0438(.A(G257), .B(new_n360), .C1(new_n331), .C2(new_n332), .ZN(new_n639));
  INV_X1    g0439(.A(G303), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n267), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n274), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n637), .A2(G179), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT84), .B1(new_n636), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n637), .A2(G179), .A3(new_n642), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n305), .A2(G116), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n490), .B2(G116), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT20), .B1(new_n634), .B2(new_n285), .ZN(new_n648));
  AND4_X1   g0448(.A1(KEYINPUT20), .A2(new_n627), .A3(new_n285), .A4(new_n629), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n645), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n637), .A2(new_n642), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G169), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n636), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n650), .A2(new_n655), .A3(KEYINPUT21), .A4(G169), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(G200), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n659), .B(new_n636), .C1(new_n277), .C2(new_n655), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n653), .A2(new_n657), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n621), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n473), .A2(new_n531), .A3(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n613), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n620), .A2(new_n613), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n577), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n576), .B1(G169), .B2(new_n584), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n578), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n613), .A4(new_n620), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n664), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(G190), .B1(new_n525), .B2(new_n526), .ZN(new_n672));
  INV_X1    g0472(.A(new_n522), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n524), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n666), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n530), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n577), .A2(new_n586), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n473), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n323), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n434), .A2(new_n285), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT11), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n436), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n442), .A2(new_n684), .A3(new_n431), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n425), .A2(G200), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT76), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n425), .A2(new_n443), .A3(G200), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n467), .ZN(new_n690));
  INV_X1    g0490(.A(new_n440), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n378), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n380), .A2(new_n354), .A3(KEYINPUT18), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n395), .B1(new_n394), .B2(new_n399), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n681), .B1(new_n696), .B2(new_n318), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n680), .A2(new_n697), .ZN(G369));
  INV_X1    g0498(.A(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n219), .A2(new_n699), .A3(new_n600), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G213), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n219), .B2(new_n600), .ZN(new_n702));
  OR3_X1    g0502(.A1(new_n701), .A2(KEYINPUT89), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT89), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n636), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n661), .B2(KEYINPUT90), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(KEYINPUT90), .B2(new_n661), .ZN(new_n711));
  INV_X1    g0511(.A(new_n676), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n709), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT91), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n531), .B1(new_n524), .B2(new_n708), .ZN(new_n717));
  INV_X1    g0517(.A(new_n530), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n708), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(G330), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n676), .A2(new_n708), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n721), .A2(new_n530), .A3(new_n523), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n530), .B2(new_n708), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n225), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n606), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n223), .A2(G50), .A3(new_n222), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n727), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT93), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n678), .B(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n671), .B1(new_n734), .B2(new_n677), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n708), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n679), .A2(new_n708), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G330), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n742));
  NOR2_X1   g0542(.A1(new_n615), .A2(G179), .ZN(new_n743));
  AND4_X1   g0543(.A1(new_n516), .A2(new_n579), .A3(new_n655), .A4(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n645), .A2(new_n519), .A3(new_n615), .A4(new_n584), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT30), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n508), .A2(new_n515), .A3(new_n615), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n643), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n584), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n744), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n708), .ZN(new_n752));
  MUX2_X1   g0552(.A(KEYINPUT31), .B(new_n742), .S(new_n752), .Z(new_n753));
  NAND3_X1  g0553(.A1(new_n662), .A2(new_n531), .A3(new_n708), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n741), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n732), .B1(new_n756), .B2(G1), .ZN(G364));
  NAND2_X1  g0557(.A1(new_n716), .A2(G330), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n329), .A2(new_n599), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G45), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G1), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n726), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n716), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n714), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n763), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n725), .A2(new_n333), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(G355), .B1(new_n628), .B2(new_n725), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n333), .A2(new_n225), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G45), .B2(new_n730), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n245), .A2(new_n254), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n220), .B1(G20), .B2(new_n320), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n770), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n219), .B1(G190), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G97), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n445), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n329), .A2(new_n277), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G107), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(G20), .A3(G190), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n333), .B1(new_n790), .B2(G87), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n784), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n219), .A2(new_n465), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(new_n445), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n277), .A3(new_n445), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n796), .A2(G58), .B1(G77), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n793), .A2(G200), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n793), .A2(KEYINPUT97), .A3(G200), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n805), .A3(G190), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n805), .A3(new_n277), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G50), .A2(new_n807), .B1(new_n809), .B2(G68), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n329), .A2(new_n277), .A3(new_n781), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  AND4_X1   g0614(.A1(new_n792), .A2(new_n801), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT98), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  INV_X1    g0617(.A(G329), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n817), .A2(new_n786), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n333), .B1(new_n640), .B2(new_n789), .C1(new_n797), .C2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G294), .C2(new_n783), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n796), .A2(G322), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT33), .B(G317), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n809), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n807), .A2(G326), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n822), .A2(new_n823), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n816), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(KEYINPUT98), .B2(new_n815), .ZN(new_n829));
  INV_X1    g0629(.A(new_n778), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n769), .B(new_n780), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT99), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n765), .A2(new_n832), .ZN(G396));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n767), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n784), .B(new_n333), .C1(new_n450), .C2(new_n789), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n209), .A2(new_n786), .B1(new_n811), .B2(new_n820), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n800), .A2(G116), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n840), .B2(new_n795), .C1(new_n640), .C2(new_n806), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n809), .A2(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n809), .A2(KEYINPUT100), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n841), .B1(G283), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n796), .A2(G143), .B1(G159), .B2(new_n800), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G150), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n847), .B2(new_n806), .C1(new_n848), .C2(new_n808), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT34), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n786), .A2(new_n207), .B1(new_n306), .B2(new_n789), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n267), .B1(new_n811), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT101), .Z(new_n854));
  AOI211_X1 g0654(.A(new_n851), .B(new_n854), .C1(G58), .C2(new_n783), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n845), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n763), .B1(G77), .B2(new_n834), .C1(new_n856), .C2(new_n830), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n463), .A2(new_n707), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n471), .A2(new_n467), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n454), .A2(new_n463), .A3(new_n466), .A4(new_n707), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n767), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n859), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n738), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n679), .A2(new_n708), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n770), .B1(new_n872), .B2(new_n755), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n755), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  INV_X1    g0676(.A(new_n544), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(G116), .A4(new_n221), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OR3_X1    g0681(.A1(new_n730), .A2(new_n266), .A3(new_n340), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n306), .A2(G68), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n304), .B(G13), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT108), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n749), .B1(new_n748), .B2(new_n584), .ZN(new_n889));
  NOR4_X1   g0689(.A1(new_n747), .A2(new_n570), .A3(new_n643), .A4(KEYINPUT30), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n886), .B(new_n888), .C1(new_n891), .C2(new_n744), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT108), .B1(new_n751), .B2(new_n887), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n742), .B1(new_n751), .B2(new_n708), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n754), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n865), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT104), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n689), .A2(new_n428), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n441), .A2(new_n708), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n440), .A2(new_n447), .A3(new_n901), .ZN(new_n904));
  OAI211_X1 g0704(.A(KEYINPUT104), .B(new_n900), .C1(new_n689), .C2(new_n428), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n904), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n415), .A2(new_n424), .A3(new_n427), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n447), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT104), .B1(new_n909), .B2(new_n900), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT105), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n897), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n267), .A2(new_n328), .A3(G20), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT7), .B1(new_n219), .B2(new_n333), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(KEYINPUT77), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n207), .B1(new_n915), .B2(new_n391), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n285), .B1(new_n916), .B2(new_n388), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT16), .B1(new_n338), .B2(new_n351), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n326), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n705), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n404), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n919), .A2(new_n920), .B1(new_n354), .B2(new_n373), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n399), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n394), .A2(new_n399), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n394), .A2(new_n920), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(new_n924), .A4(new_n374), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n923), .A2(new_n935), .A3(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT38), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT79), .B1(new_n693), .B2(new_n694), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n401), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n921), .B1(new_n939), .B2(new_n378), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n363), .A2(new_n277), .A3(new_n368), .ZN(new_n941));
  AOI21_X1  g0741(.A(G200), .B1(new_n363), .B2(new_n368), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n394), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n346), .A2(new_n353), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n945), .A2(new_n326), .B1(new_n397), .B2(new_n398), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n947), .A2(KEYINPUT106), .A3(new_n924), .A4(new_n930), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n931), .A2(new_n932), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n927), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n937), .B1(new_n940), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n936), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT40), .B1(new_n912), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n929), .A2(new_n930), .A3(new_n374), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n948), .A2(new_n949), .B1(KEYINPUT37), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n930), .B1(new_n378), .B2(new_n695), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n937), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n954), .B1(new_n936), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n953), .B1(new_n912), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n473), .A2(new_n896), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(G330), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(KEYINPUT109), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(KEYINPUT109), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n940), .A2(new_n950), .A3(new_n937), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n955), .A2(KEYINPUT37), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n933), .B2(new_n934), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n378), .A2(new_n695), .ZN(new_n970));
  INV_X1    g0770(.A(new_n930), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT38), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n966), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n691), .A2(new_n708), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n936), .A2(new_n951), .A3(KEYINPUT39), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT107), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n695), .A2(new_n920), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n464), .A2(new_n466), .A3(new_n708), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n906), .A2(new_n911), .B1(new_n870), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n980), .B1(new_n982), .B2(new_n952), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n978), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n979), .B1(new_n978), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n473), .B1(new_n737), .B2(new_n739), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n697), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n986), .B(new_n988), .Z(new_n989));
  OAI22_X1  g0789(.A1(new_n965), .A2(new_n989), .B1(new_n304), .B2(new_n760), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n965), .A2(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n885), .B1(new_n990), .B2(new_n991), .ZN(G367));
  NAND2_X1  g0792(.A1(new_n774), .A2(new_n237), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n778), .B(new_n768), .C1(new_n725), .C2(new_n456), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n770), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n768), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n618), .A2(new_n601), .A3(new_n619), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n675), .B1(new_n998), .B2(new_n708), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n664), .A2(new_n997), .A3(new_n707), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n807), .A2(G143), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n811), .A2(new_n847), .B1(new_n339), .B2(new_n789), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT113), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n783), .A2(G68), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n333), .B1(new_n787), .B2(G77), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n796), .A2(G150), .B1(G50), .B2(new_n800), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G159), .C2(new_n844), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n796), .A2(G303), .B1(G283), .B2(new_n800), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n787), .A2(G97), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n450), .B2(new_n782), .C1(new_n1014), .C2(new_n811), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n790), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT46), .B1(new_n790), .B2(G116), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1015), .A2(new_n267), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1012), .B(new_n1018), .C1(new_n820), .C2(new_n806), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G294), .B2(new_n844), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1011), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT47), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n995), .B1(new_n996), .B2(new_n1001), .C1(new_n1022), .C2(new_n830), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n720), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n678), .B(KEYINPUT93), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n578), .B2(new_n708), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n577), .A2(new_n708), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT110), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(KEYINPUT45), .A3(new_n723), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n723), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n723), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT44), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT44), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1029), .B2(new_n723), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1030), .A2(new_n1033), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT111), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1024), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1033), .A2(new_n1030), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(KEYINPUT111), .A3(new_n720), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n758), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n716), .A2(KEYINPUT112), .A3(G330), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n722), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n721), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n719), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n1052), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1046), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n756), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n726), .B(KEYINPUT41), .Z(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n762), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1034), .A2(KEYINPUT42), .A3(new_n1050), .ZN(new_n1062));
  OAI21_X1  g0862(.A(KEYINPUT42), .B1(new_n1034), .B2(new_n1050), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT43), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1001), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n577), .B1(new_n1034), .B2(new_n718), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n708), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n1063), .A3(new_n1062), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1066), .A2(new_n1065), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1073), .A2(new_n1024), .A3(new_n1029), .A4(new_n1069), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1023), .B1(new_n1061), .B2(new_n1078), .ZN(G387));
  NAND2_X1  g0879(.A1(new_n1056), .A2(new_n756), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n756), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n726), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n719), .A2(new_n996), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n728), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(new_n771), .B1(new_n450), .B2(new_n725), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n234), .A2(new_n254), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n295), .A2(new_n306), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT50), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n728), .B(new_n254), .C1(new_n207), .C2(new_n266), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n774), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1086), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n779), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n763), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n797), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n809), .A2(new_n295), .B1(G68), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT114), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n782), .A2(new_n455), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n811), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(G150), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n790), .A2(G77), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1100), .A2(new_n267), .A3(new_n1013), .A4(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n796), .B2(G50), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1097), .B(new_n1103), .C1(new_n812), .C2(new_n806), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n267), .B1(new_n1099), .B2(G326), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n782), .A2(new_n817), .B1(new_n840), .B2(new_n789), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G303), .A2(new_n800), .B1(new_n796), .B2(G317), .ZN(new_n1107));
  INV_X1    g0907(.A(G322), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n844), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n806), .C1(new_n1109), .C2(new_n820), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT48), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1111), .B2(new_n1110), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT49), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1105), .B1(new_n628), .B2(new_n786), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1104), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1084), .B(new_n1094), .C1(new_n1117), .C2(new_n778), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1056), .B2(new_n762), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1083), .A2(new_n1119), .ZN(G393));
  XNOR2_X1  g0920(.A(new_n1044), .B(new_n720), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n727), .B1(new_n1056), .B2(new_n756), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n762), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1041), .A2(new_n1045), .A3(new_n726), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1081), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1034), .A2(new_n768), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n774), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n242), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n779), .B1(new_n550), .B2(new_n225), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n763), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n795), .A2(new_n812), .B1(new_n848), .B2(new_n806), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n844), .A2(G50), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n782), .A2(new_n266), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G143), .B2(new_n1099), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n333), .B1(new_n790), .B2(G68), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n209), .C2(new_n786), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n295), .B2(new_n800), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1135), .A2(new_n1136), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n782), .A2(new_n628), .B1(new_n811), .B2(new_n1108), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n788), .B(new_n333), .C1(new_n817), .C2(new_n789), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(G294), .C2(new_n1095), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1109), .B2(new_n640), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n795), .A2(new_n820), .B1(new_n1014), .B2(new_n806), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1143), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1131), .B1(new_n1151), .B2(new_n778), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1125), .A2(new_n1126), .B1(new_n1127), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1123), .A2(new_n1153), .ZN(G390));
  INV_X1    g0954(.A(G125), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n306), .A2(new_n786), .B1(new_n811), .B2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1157));
  AND3_X1   g0957(.A1(new_n790), .A2(G150), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n790), .B2(G150), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .A4(new_n333), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n795), .B2(new_n852), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n800), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1162), .A2(new_n1163), .B1(new_n812), .B2(new_n782), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n844), .B2(G137), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT118), .Z(new_n1166));
  AOI211_X1 g0966(.A(new_n1161), .B(new_n1166), .C1(G128), .C2(new_n807), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n333), .B1(new_n209), .B2(new_n789), .C1(new_n786), .C2(new_n207), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n782), .A2(new_n266), .B1(new_n811), .B2(new_n840), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n796), .C2(G116), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n550), .B2(new_n1162), .C1(new_n817), .C2(new_n806), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G107), .B2(new_n844), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n778), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n763), .C1(new_n295), .C2(new_n834), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n974), .A2(new_n977), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n766), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n897), .A2(new_n741), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n911), .A2(new_n906), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n870), .A2(new_n981), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n974), .A2(new_n977), .B1(new_n1181), .B2(new_n975), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n981), .B1(new_n736), .B2(new_n868), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1178), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n976), .B1(new_n936), .B2(new_n958), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1181), .A2(new_n975), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1175), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n755), .A2(new_n1178), .A3(new_n865), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1187), .A2(KEYINPUT117), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT117), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n1179), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1176), .B1(new_n1197), .B2(new_n762), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1178), .B1(new_n755), .B2(new_n865), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1180), .B1(new_n1179), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1183), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1191), .B(new_n1201), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n473), .A2(G330), .A3(new_n896), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n987), .A2(new_n1204), .A3(new_n697), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n726), .B1(new_n1197), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1198), .B1(new_n1209), .B2(new_n1210), .ZN(G378));
  AOI21_X1  g1011(.A(new_n705), .B1(new_n303), .B2(new_n310), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n324), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n681), .B1(new_n314), .B2(new_n317), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1212), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n681), .B(new_n1212), .C1(new_n314), .C2(new_n317), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n766), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n763), .B1(G50), .B2(new_n834), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n783), .A2(G150), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n847), .B2(new_n797), .C1(new_n789), .C2(new_n1163), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n796), .B2(G128), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n1155), .B2(new_n806), .C1(new_n852), .C2(new_n808), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n282), .B(new_n253), .C1(new_n786), .C2(new_n812), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G124), .B2(new_n1099), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1006), .A2(new_n253), .A3(new_n333), .A4(new_n1101), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n786), .A2(new_n339), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G283), .B2(new_n1099), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n455), .B2(new_n797), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1235), .B(new_n1238), .C1(new_n796), .C2(G107), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n550), .B2(new_n808), .C1(new_n628), .C2(new_n806), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G50), .B1(new_n282), .B2(new_n253), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n267), .B2(G41), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT120), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1234), .A2(new_n1242), .A3(new_n1243), .A4(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1225), .B1(new_n1247), .B2(new_n778), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1224), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT40), .B1(new_n967), .B2(new_n973), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n896), .A2(new_n865), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1178), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(G330), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1254), .A2(new_n953), .A3(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n936), .A2(new_n951), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n954), .B1(new_n1257), .B2(new_n1253), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n741), .B1(new_n912), .B2(new_n959), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1223), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1256), .A2(new_n1260), .B1(new_n984), .B2(new_n985), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT121), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n978), .A2(new_n983), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT107), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1255), .B1(new_n1254), .B2(new_n953), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n978), .A2(new_n983), .A3(new_n979), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1258), .A2(new_n1259), .A3(new_n1223), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n986), .A2(KEYINPUT121), .A3(new_n1267), .A4(new_n1265), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1250), .B1(new_n1271), .B2(new_n762), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1273));
  AOI211_X1 g1073(.A(KEYINPUT117), .B(new_n1273), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1195), .B1(new_n1194), .B2(new_n1179), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1192), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1206), .B1(new_n1276), .B2(new_n1207), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1210), .A2(new_n1205), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT57), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1261), .B2(new_n1268), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n726), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1272), .B1(new_n1278), .B2(new_n1283), .ZN(G375));
  NAND3_X1  g1084(.A1(new_n1200), .A2(new_n1205), .A3(new_n1202), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT122), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1200), .A2(KEYINPUT122), .A3(new_n1205), .A4(new_n1202), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1060), .A3(new_n1207), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1203), .A2(new_n762), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n763), .B1(G68), .B2(new_n834), .ZN(new_n1292));
  OAI221_X1 g1092(.A(new_n333), .B1(new_n550), .B2(new_n789), .C1(new_n786), .C2(new_n266), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n782), .A2(new_n455), .B1(new_n811), .B2(new_n640), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n1293), .B(new_n1294), .C1(new_n796), .C2(G283), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n1295), .B1(new_n450), .B2(new_n1162), .C1(new_n840), .C2(new_n806), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1109), .A2(new_n628), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1109), .A2(new_n1163), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n267), .B1(new_n812), .B2(new_n789), .C1(new_n786), .C2(new_n339), .ZN(new_n1299));
  INV_X1    g1099(.A(G128), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n797), .A2(new_n848), .B1(new_n1300), .B2(new_n811), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1299), .B(new_n1301), .C1(G50), .C2(new_n783), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1302), .B1(new_n852), .B2(new_n806), .C1(new_n847), .C2(new_n795), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n1296), .A2(new_n1297), .B1(new_n1298), .B2(new_n1303), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1304), .A2(KEYINPUT123), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n830), .B1(new_n1304), .B2(KEYINPUT123), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1292), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1178), .B2(new_n767), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1291), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(new_n1310), .ZN(G381));
  INV_X1    g1111(.A(G396), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1083), .A2(new_n1312), .A3(new_n1119), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(G384), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(KEYINPUT124), .ZN(new_n1315));
  INV_X1    g1115(.A(G378), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n762), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1249), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n727), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1270), .B(new_n1269), .C1(new_n1210), .C2(new_n1205), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1280), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(G387), .A2(G381), .A3(G390), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1315), .A2(new_n1316), .A3(new_n1323), .A4(new_n1324), .ZN(G407));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n706), .A3(new_n1316), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G407), .A2(G213), .A3(new_n1326), .ZN(G409));
  INV_X1    g1127(.A(G213), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1328), .A2(G343), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(G2897), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1207), .A2(KEYINPUT60), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT60), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n726), .B1(new_n1285), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1332), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G384), .B1(new_n1336), .B2(new_n1310), .ZN(new_n1337));
  AOI211_X1 g1137(.A(new_n875), .B(new_n1309), .C1(new_n1332), .C2(new_n1335), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1330), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1334), .B1(new_n1289), .B2(new_n1331), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n875), .B1(new_n1340), .B2(new_n1309), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1336), .A2(G384), .A3(new_n1310), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1341), .A2(G2897), .A3(new_n1342), .A4(new_n1329), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1344));
  OAI211_X1 g1144(.A(G378), .B(new_n1272), .C1(new_n1278), .C2(new_n1283), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1261), .A2(new_n1268), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1250), .B1(new_n1346), .B2(new_n762), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1347), .B1(new_n1321), .B2(new_n1059), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1316), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1329), .B1(new_n1345), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT125), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1344), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1271), .A2(new_n1277), .A3(new_n1060), .ZN(new_n1353));
  AOI21_X1  g1153(.A(G378), .B1(new_n1353), .B2(new_n1347), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(G378), .B2(new_n1323), .ZN(new_n1355));
  OAI21_X1  g1155(.A(KEYINPUT125), .B1(new_n1355), .B2(new_n1329), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1352), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT61), .ZN(new_n1358));
  AOI22_X1  g1158(.A1(new_n1041), .A2(new_n1045), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1060), .B1(new_n1359), .B2(new_n1081), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1078), .B1(new_n1318), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1023), .ZN(new_n1362));
  OAI21_X1  g1162(.A(KEYINPUT126), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT126), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1364), .B(new_n1023), .C1(new_n1061), .C2(new_n1078), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1127), .A2(new_n1152), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1366), .B1(new_n1080), .B2(new_n1124), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1318), .B1(new_n1126), .B2(new_n727), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1367), .B1(new_n1368), .B2(new_n1121), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1083), .A2(new_n1312), .A3(new_n1119), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1312), .B1(new_n1083), .B2(new_n1119), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1369), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(G393), .A2(G396), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1373), .A2(G390), .A3(new_n1313), .ZN(new_n1374));
  AND4_X1   g1174(.A1(new_n1363), .A2(new_n1365), .A3(new_n1372), .A4(new_n1374), .ZN(new_n1375));
  AOI22_X1  g1175(.A1(new_n1363), .A2(new_n1365), .B1(new_n1372), .B2(new_n1374), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1358), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1345), .A2(new_n1349), .ZN(new_n1378));
  INV_X1    g1178(.A(new_n1329), .ZN(new_n1379));
  NOR2_X1   g1179(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1378), .A2(new_n1379), .A3(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT63), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1377), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1350), .A2(KEYINPUT63), .A3(new_n1380), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1357), .A2(new_n1383), .A3(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT62), .ZN(new_n1386));
  AND3_X1   g1186(.A1(new_n1350), .A2(new_n1386), .A3(new_n1380), .ZN(new_n1387));
  OAI21_X1  g1187(.A(new_n1358), .B1(new_n1350), .B2(new_n1344), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1386), .B1(new_n1350), .B2(new_n1380), .ZN(new_n1389));
  NOR3_X1   g1189(.A1(new_n1387), .A2(new_n1388), .A3(new_n1389), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1391));
  INV_X1    g1191(.A(new_n1391), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n1385), .B1(new_n1390), .B2(new_n1392), .ZN(G405));
  NOR2_X1   g1193(.A1(new_n1323), .A2(G378), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1345), .ZN(new_n1395));
  OR3_X1    g1195(.A1(new_n1394), .A2(new_n1395), .A3(new_n1380), .ZN(new_n1396));
  OAI21_X1  g1196(.A(new_n1380), .B1(new_n1394), .B2(new_n1395), .ZN(new_n1397));
  AND3_X1   g1197(.A1(new_n1396), .A2(new_n1391), .A3(new_n1397), .ZN(new_n1398));
  AOI21_X1  g1198(.A(new_n1391), .B1(new_n1396), .B2(new_n1397), .ZN(new_n1399));
  NOR2_X1   g1199(.A1(new_n1398), .A2(new_n1399), .ZN(G402));
endmodule


