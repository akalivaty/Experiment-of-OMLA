

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577;

  NOR2_X1 U321 ( .A1(n445), .A2(n435), .ZN(n557) );
  XNOR2_X1 U322 ( .A(KEYINPUT48), .B(n402), .ZN(n535) );
  XNOR2_X1 U323 ( .A(n355), .B(n354), .ZN(n356) );
  NOR2_X1 U324 ( .A1(n536), .A2(n416), .ZN(n563) );
  XNOR2_X1 U325 ( .A(n357), .B(n356), .ZN(n358) );
  INV_X1 U326 ( .A(G190GAT), .ZN(n436) );
  XNOR2_X1 U327 ( .A(n344), .B(n343), .ZN(n564) );
  XNOR2_X1 U328 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U329 ( .A(n439), .B(n438), .ZN(G1351GAT) );
  XNOR2_X1 U330 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n289) );
  XNOR2_X1 U331 ( .A(n289), .B(KEYINPUT78), .ZN(n290) );
  XOR2_X1 U332 ( .A(n290), .B(KEYINPUT17), .Z(n292) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n410) );
  XOR2_X1 U335 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n294) );
  XNOR2_X1 U336 ( .A(G15GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(n295), .B(G190GAT), .Z(n297) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n389) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(n389), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U342 ( .A(KEYINPUT80), .B(G176GAT), .Z(n299) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U345 ( .A(n301), .B(n300), .Z(n307) );
  XNOR2_X1 U346 ( .A(G127GAT), .B(KEYINPUT75), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n302), .B(KEYINPUT0), .ZN(n303) );
  XOR2_X1 U348 ( .A(n303), .B(KEYINPUT76), .Z(n305) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(G134GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n325) );
  XNOR2_X1 U351 ( .A(n325), .B(KEYINPUT77), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n410), .B(n308), .ZN(n445) );
  XNOR2_X1 U354 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n434) );
  XOR2_X1 U355 ( .A(KEYINPUT1), .B(G120GAT), .Z(n310) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(G1GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n312) );
  XNOR2_X1 U359 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT83), .B(KEYINPUT6), .Z(n316) );
  NAND2_X1 U363 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U365 ( .A(G57GAT), .B(n317), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G162GAT), .Z(n322) );
  XNOR2_X1 U368 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n320), .B(KEYINPUT3), .ZN(n429) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(n429), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U372 ( .A(n324), .B(n323), .Z(n327) );
  XNOR2_X1 U373 ( .A(n325), .B(G148GAT), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n536) );
  XOR2_X1 U375 ( .A(G197GAT), .B(G50GAT), .Z(n329) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(G36GAT), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U378 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n331) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n344) );
  XOR2_X1 U382 ( .A(G141GAT), .B(G22GAT), .Z(n417) );
  XOR2_X1 U383 ( .A(KEYINPUT68), .B(G8GAT), .Z(n335) );
  XNOR2_X1 U384 ( .A(G15GAT), .B(G1GAT), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n372) );
  XOR2_X1 U386 ( .A(n417), .B(n372), .Z(n337) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(n338), .B(KEYINPUT65), .Z(n342) );
  XOR2_X1 U390 ( .A(G29GAT), .B(G43GAT), .Z(n340) );
  XNOR2_X1 U391 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n347) );
  XNOR2_X1 U393 ( .A(n347), .B(KEYINPUT30), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U395 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n346) );
  XNOR2_X1 U396 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U398 ( .A(G99GAT), .B(G85GAT), .Z(n388) );
  XNOR2_X1 U399 ( .A(n347), .B(n388), .ZN(n349) );
  AND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n357) );
  XNOR2_X1 U402 ( .A(G50GAT), .B(KEYINPUT70), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n350), .B(G162GAT), .ZN(n422) );
  XNOR2_X1 U404 ( .A(G36GAT), .B(G190GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n351), .B(G218GAT), .ZN(n403) );
  XNOR2_X1 U406 ( .A(n422), .B(n403), .ZN(n355) );
  XOR2_X1 U407 ( .A(G92GAT), .B(KEYINPUT64), .Z(n353) );
  XNOR2_X1 U408 ( .A(G134GAT), .B(G106GAT), .ZN(n352) );
  XOR2_X1 U409 ( .A(n353), .B(n352), .Z(n354) );
  XOR2_X1 U410 ( .A(n359), .B(n358), .Z(n547) );
  XOR2_X1 U411 ( .A(KEYINPUT36), .B(n547), .Z(n574) );
  XOR2_X1 U412 ( .A(G64GAT), .B(G71GAT), .Z(n361) );
  XNOR2_X1 U413 ( .A(G183GAT), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n376) );
  XOR2_X1 U415 ( .A(G211GAT), .B(G155GAT), .Z(n363) );
  XNOR2_X1 U416 ( .A(G22GAT), .B(G78GAT), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n368) );
  XNOR2_X1 U418 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n364), .B(KEYINPUT69), .ZN(n386) );
  XOR2_X1 U420 ( .A(KEYINPUT12), .B(n386), .Z(n366) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n374) );
  XOR2_X1 U424 ( .A(KEYINPUT73), .B(KEYINPUT15), .Z(n370) );
  XNOR2_X1 U425 ( .A(KEYINPUT14), .B(KEYINPUT72), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n472) );
  NOR2_X1 U430 ( .A1(n574), .A2(n472), .ZN(n377) );
  XNOR2_X1 U431 ( .A(KEYINPUT45), .B(n377), .ZN(n392) );
  XOR2_X1 U432 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n379) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(n380), .B(KEYINPUT31), .Z(n385) );
  XNOR2_X1 U436 ( .A(G106GAT), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n381), .B(G148GAT), .ZN(n430) );
  XOR2_X1 U438 ( .A(G64GAT), .B(G92GAT), .Z(n383) );
  XNOR2_X1 U439 ( .A(G176GAT), .B(G204GAT), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n406) );
  XNOR2_X1 U441 ( .A(n430), .B(n406), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U443 ( .A(n387), .B(n386), .Z(n391) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n567) );
  NAND2_X1 U446 ( .A1(n392), .A2(n567), .ZN(n393) );
  NOR2_X1 U447 ( .A1(n564), .A2(n393), .ZN(n394) );
  XOR2_X1 U448 ( .A(n394), .B(KEYINPUT109), .Z(n401) );
  XNOR2_X1 U449 ( .A(KEYINPUT41), .B(n567), .ZN(n554) );
  NAND2_X1 U450 ( .A1(n564), .A2(n554), .ZN(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U453 ( .A1(n397), .A2(n472), .ZN(n398) );
  NOR2_X1 U454 ( .A1(n547), .A2(n398), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT47), .B(n399), .Z(n400) );
  NOR2_X1 U456 ( .A1(n401), .A2(n400), .ZN(n402) );
  XOR2_X1 U457 ( .A(n403), .B(G8GAT), .Z(n405) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U460 ( .A(n407), .B(n406), .Z(n412) );
  XOR2_X1 U461 ( .A(G211GAT), .B(KEYINPUT21), .Z(n409) );
  XNOR2_X1 U462 ( .A(G197GAT), .B(KEYINPUT81), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n410), .B(n418), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n507) );
  XOR2_X1 U466 ( .A(KEYINPUT120), .B(n507), .Z(n413) );
  NOR2_X1 U467 ( .A1(n535), .A2(n413), .ZN(n415) );
  INV_X1 U468 ( .A(KEYINPUT54), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U470 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U473 ( .A(n421), .B(G204GAT), .Z(n424) );
  XNOR2_X1 U474 ( .A(n422), .B(KEYINPUT22), .ZN(n423) );
  XNOR2_X1 U475 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U476 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n426) );
  XNOR2_X1 U477 ( .A(G218GAT), .B(KEYINPUT82), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U479 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U480 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U481 ( .A(n432), .B(n431), .ZN(n449) );
  NAND2_X1 U482 ( .A1(n563), .A2(n449), .ZN(n433) );
  XNOR2_X1 U483 ( .A(n434), .B(n433), .ZN(n435) );
  NAND2_X1 U484 ( .A1(n557), .A2(n547), .ZN(n439) );
  XOR2_X1 U485 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n437) );
  XOR2_X1 U486 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n462) );
  XOR2_X1 U487 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n441) );
  OR2_X1 U488 ( .A1(n472), .A2(n547), .ZN(n440) );
  XNOR2_X1 U489 ( .A(n441), .B(n440), .ZN(n459) );
  XOR2_X1 U490 ( .A(n449), .B(KEYINPUT28), .Z(n511) );
  XOR2_X1 U491 ( .A(n507), .B(KEYINPUT86), .Z(n442) );
  XNOR2_X1 U492 ( .A(KEYINPUT27), .B(n442), .ZN(n452) );
  NOR2_X1 U493 ( .A1(n511), .A2(n452), .ZN(n443) );
  NAND2_X1 U494 ( .A1(n536), .A2(n443), .ZN(n517) );
  XNOR2_X1 U495 ( .A(n517), .B(KEYINPUT87), .ZN(n444) );
  NAND2_X1 U496 ( .A1(n444), .A2(n445), .ZN(n458) );
  INV_X1 U497 ( .A(n445), .ZN(n518) );
  NAND2_X1 U498 ( .A1(n507), .A2(n518), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n446), .A2(n449), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n447), .B(KEYINPUT25), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n448), .B(KEYINPUT89), .ZN(n454) );
  XNOR2_X1 U502 ( .A(KEYINPUT26), .B(KEYINPUT88), .ZN(n451) );
  NOR2_X1 U503 ( .A1(n518), .A2(n449), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n562) );
  INV_X1 U505 ( .A(n452), .ZN(n453) );
  NAND2_X1 U506 ( .A1(n562), .A2(n453), .ZN(n534) );
  NAND2_X1 U507 ( .A1(n454), .A2(n534), .ZN(n456) );
  INV_X1 U508 ( .A(n536), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n456), .A2(n455), .ZN(n457) );
  NAND2_X1 U510 ( .A1(n458), .A2(n457), .ZN(n474) );
  NAND2_X1 U511 ( .A1(n459), .A2(n474), .ZN(n491) );
  NAND2_X1 U512 ( .A1(n564), .A2(n567), .ZN(n477) );
  NOR2_X1 U513 ( .A1(n491), .A2(n477), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT90), .ZN(n469) );
  NAND2_X1 U515 ( .A1(n536), .A2(n469), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U517 ( .A(G1GAT), .B(n463), .ZN(G1324GAT) );
  NAND2_X1 U518 ( .A1(n469), .A2(n507), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U520 ( .A(KEYINPUT35), .B(KEYINPUT93), .Z(n466) );
  NAND2_X1 U521 ( .A1(n518), .A2(n469), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n468) );
  XOR2_X1 U523 ( .A(G15GAT), .B(KEYINPUT92), .Z(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(G1326GAT) );
  NAND2_X1 U525 ( .A1(n469), .A2(n511), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT94), .ZN(n471) );
  XNOR2_X1 U527 ( .A(G22GAT), .B(n471), .ZN(G1327GAT) );
  XOR2_X1 U528 ( .A(G29GAT), .B(KEYINPUT39), .Z(n480) );
  INV_X1 U529 ( .A(n472), .ZN(n570) );
  NOR2_X1 U530 ( .A1(n570), .A2(n574), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT37), .B(n475), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT95), .B(n476), .ZN(n504) );
  NOR2_X1 U534 ( .A1(n477), .A2(n504), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT38), .ZN(n486) );
  NAND2_X1 U536 ( .A1(n536), .A2(n486), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(G1328GAT) );
  NAND2_X1 U538 ( .A1(n486), .A2(n507), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G36GAT), .B(n482), .ZN(G1329GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT40), .B(KEYINPUT97), .Z(n484) );
  NAND2_X1 U542 ( .A1(n518), .A2(n486), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G43GAT), .B(n485), .ZN(G1330GAT) );
  NAND2_X1 U545 ( .A1(n486), .A2(n511), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U547 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT99), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT98), .B(n489), .Z(n493) );
  INV_X1 U550 ( .A(n564), .ZN(n490) );
  NAND2_X1 U551 ( .A1(n490), .A2(n554), .ZN(n503) );
  NOR2_X1 U552 ( .A1(n491), .A2(n503), .ZN(n498) );
  NAND2_X1 U553 ( .A1(n498), .A2(n536), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1332GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n507), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(KEYINPUT100), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G64GAT), .B(n495), .ZN(G1333GAT) );
  XOR2_X1 U558 ( .A(G71GAT), .B(KEYINPUT101), .Z(n497) );
  NAND2_X1 U559 ( .A1(n498), .A2(n518), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1334GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n500) );
  NAND2_X1 U562 ( .A1(n498), .A2(n511), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n502) );
  XOR2_X1 U564 ( .A(G78GAT), .B(KEYINPUT103), .Z(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  XNOR2_X1 U566 ( .A(G85GAT), .B(KEYINPUT104), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n504), .A2(n503), .ZN(n512) );
  NAND2_X1 U568 ( .A1(n536), .A2(n512), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1336GAT) );
  XOR2_X1 U570 ( .A(G92GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U571 ( .A1(n512), .A2(n507), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1337GAT) );
  NAND2_X1 U573 ( .A1(n512), .A2(n518), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U575 ( .A(G106GAT), .B(KEYINPUT106), .ZN(n516) );
  XOR2_X1 U576 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n514) );
  NAND2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1339GAT) );
  XOR2_X1 U580 ( .A(G113GAT), .B(KEYINPUT111), .Z(n522) );
  NOR2_X1 U581 ( .A1(n535), .A2(n517), .ZN(n519) );
  NAND2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(n520), .Z(n529) );
  NAND2_X1 U584 ( .A1(n564), .A2(n529), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(G120GAT), .B(KEYINPUT49), .Z(n524) );
  NAND2_X1 U587 ( .A1(n529), .A2(n554), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1341GAT) );
  XNOR2_X1 U589 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n528) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n526) );
  NAND2_X1 U591 ( .A1(n570), .A2(n529), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1342GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U595 ( .A1(n547), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT114), .Z(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1343GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(n538), .Z(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n564), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n541) );
  NAND2_X1 U605 ( .A1(n546), .A2(n554), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT53), .Z(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n546), .A2(n570), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(KEYINPUT118), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G155GAT), .B(n545), .ZN(G1346GAT) );
  XOR2_X1 U612 ( .A(G162GAT), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n557), .A2(n564), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT122), .B(n553), .Z(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n570), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n560) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(n561), .Z(n566) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n573) );
  INV_X1 U630 ( .A(n573), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n571), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .Z(n569) );
  OR2_X1 U634 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1353GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(n577), .ZN(G1355GAT) );
endmodule

