

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U555 ( .A1(n629), .A2(n733), .ZN(n699) );
  XNOR2_X1 U556 ( .A(n661), .B(KEYINPUT15), .ZN(n662) );
  AND2_X1 U557 ( .A1(n733), .A2(G2072), .ZN(n558) );
  AND2_X1 U558 ( .A1(n551), .A2(n549), .ZN(n548) );
  INV_X1 U559 ( .A(n699), .ZN(n680) );
  OR2_X1 U560 ( .A1(n695), .A2(n694), .ZN(n696) );
  AND2_X1 U561 ( .A1(n724), .A2(n723), .ZN(n541) );
  AND2_X1 U562 ( .A1(n728), .A2(n539), .ZN(n538) );
  INV_X1 U563 ( .A(KEYINPUT33), .ZN(n539) );
  AND2_X1 U564 ( .A1(n563), .A2(n762), .ZN(n763) );
  NOR2_X1 U565 ( .A1(n533), .A2(n532), .ZN(n531) );
  INV_X1 U566 ( .A(n763), .ZN(n533) );
  NOR2_X1 U567 ( .A1(n763), .A2(KEYINPUT99), .ZN(n529) );
  INV_X1 U568 ( .A(KEYINPUT99), .ZN(n532) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n628) );
  NAND2_X1 U570 ( .A1(n626), .A2(n625), .ZN(n537) );
  INV_X1 U571 ( .A(KEYINPUT85), .ZN(n536) );
  AND2_X1 U572 ( .A1(n561), .A2(n566), .ZN(n560) );
  XNOR2_X1 U573 ( .A(n562), .B(KEYINPUT66), .ZN(n561) );
  XNOR2_X1 U574 ( .A(n559), .B(n630), .ZN(n632) );
  NAND2_X1 U575 ( .A1(n546), .A2(n545), .ZN(n544) );
  AND2_X1 U576 ( .A1(G286), .A2(n697), .ZN(n552) );
  AND2_X1 U577 ( .A1(n550), .A2(n703), .ZN(n549) );
  OR2_X1 U578 ( .A1(G286), .A2(n697), .ZN(n550) );
  NOR2_X1 U579 ( .A1(n706), .A2(n705), .ZN(n709) );
  INV_X1 U580 ( .A(n998), .ZN(n557) );
  NAND2_X1 U581 ( .A1(n543), .A2(n565), .ZN(n542) );
  INV_X1 U582 ( .A(G2104), .ZN(n543) );
  AND2_X1 U583 ( .A1(n530), .A2(n528), .ZN(n527) );
  NOR2_X1 U584 ( .A1(n529), .A2(n524), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n526), .A2(n532), .ZN(n525) );
  XNOR2_X1 U586 ( .A(n537), .B(n536), .ZN(n535) );
  NOR2_X1 U587 ( .A1(n569), .A2(n568), .ZN(G160) );
  NAND2_X1 U588 ( .A1(n521), .A2(n560), .ZN(n569) );
  NOR2_X1 U589 ( .A1(n627), .A2(n535), .ZN(G164) );
  XOR2_X1 U590 ( .A(n564), .B(KEYINPUT23), .Z(n521) );
  AND2_X1 U591 ( .A1(n555), .A2(n721), .ZN(n522) );
  NAND2_X1 U592 ( .A1(n540), .A2(n538), .ZN(n523) );
  INV_X1 U593 ( .A(n662), .ZN(n545) );
  AND2_X1 U594 ( .A1(n994), .A2(n774), .ZN(n524) );
  INV_X1 U595 ( .A(n696), .ZN(n705) );
  NAND2_X1 U596 ( .A1(n764), .A2(n531), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n527), .A2(n525), .ZN(n534) );
  INV_X1 U598 ( .A(n764), .ZN(n526) );
  NAND2_X1 U599 ( .A1(n534), .A2(n776), .ZN(n777) );
  NAND2_X1 U600 ( .A1(n725), .A2(n541), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n704), .B(KEYINPUT32), .ZN(n725) );
  XNOR2_X2 U602 ( .A(n542), .B(KEYINPUT17), .ZN(n881) );
  NAND2_X1 U603 ( .A1(n673), .A2(n544), .ZN(n676) );
  NAND2_X1 U604 ( .A1(n666), .A2(n653), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n642), .B(n641), .ZN(n666) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n705), .A2(KEYINPUT95), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n696), .A2(n552), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n553), .A2(G8), .ZN(n704) );
  NAND2_X1 U610 ( .A1(n522), .A2(n554), .ZN(n764) );
  NAND2_X1 U611 ( .A1(n716), .A2(n698), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n523), .A2(n556), .ZN(n555) );
  NOR2_X1 U613 ( .A1(n732), .A2(n557), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n629), .A2(n558), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n881), .A2(G137), .ZN(n562) );
  NOR2_X1 U616 ( .A1(n699), .A2(n921), .ZN(n642) );
  OR2_X1 U617 ( .A1(n761), .A2(n1015), .ZN(n563) );
  AND2_X1 U618 ( .A1(n663), .A2(n652), .ZN(n653) );
  XNOR2_X1 U619 ( .A(n686), .B(KEYINPUT93), .ZN(n687) );
  XNOR2_X1 U620 ( .A(n688), .B(n687), .ZN(n689) );
  INV_X1 U621 ( .A(KEYINPUT95), .ZN(n697) );
  AND2_X1 U622 ( .A1(n565), .A2(G2104), .ZN(n882) );
  NOR2_X2 U623 ( .A1(G2104), .A2(n565), .ZN(n886) );
  NOR2_X1 U624 ( .A1(n612), .A2(G651), .ZN(n820) );
  INV_X1 U625 ( .A(G2105), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G101), .A2(n882), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n886), .A2(G125), .ZN(n566) );
  AND2_X1 U628 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U629 ( .A1(G113), .A2(n885), .ZN(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT65), .B(n567), .ZN(n568) );
  INV_X1 U631 ( .A(G651), .ZN(n573) );
  NOR2_X1 U632 ( .A1(G543), .A2(n573), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT1), .B(n570), .Z(n815) );
  NAND2_X1 U634 ( .A1(G64), .A2(n815), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT0), .B(G543), .Z(n612) );
  NAND2_X1 U636 ( .A1(G52), .A2(n820), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n578) );
  NOR2_X1 U638 ( .A1(G543), .A2(G651), .ZN(n816) );
  NAND2_X1 U639 ( .A1(G90), .A2(n816), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n612), .A2(n573), .ZN(n819) );
  NAND2_X1 U641 ( .A1(G77), .A2(n819), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT67), .B(n579), .Z(G171) );
  INV_X1 U646 ( .A(G171), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G63), .A2(n815), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G51), .A2(n820), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT6), .B(n582), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n816), .A2(G89), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT4), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G76), .A2(n819), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT5), .B(n586), .Z(n587) );
  XNOR2_X1 U656 ( .A(KEYINPUT72), .B(n587), .ZN(n588) );
  NOR2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U658 ( .A(KEYINPUT7), .B(KEYINPUT73), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n591), .B(n590), .ZN(G168) );
  XOR2_X1 U660 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U661 ( .A1(n819), .A2(G75), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT79), .B(n592), .Z(n594) );
  NAND2_X1 U663 ( .A1(n816), .A2(G88), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U665 ( .A(KEYINPUT80), .B(n595), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G50), .A2(n820), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(KEYINPUT78), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n815), .A2(G62), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G166) );
  INV_X1 U671 ( .A(G166), .ZN(G303) );
  NAND2_X1 U672 ( .A1(G61), .A2(n815), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G86), .A2(n816), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G73), .A2(n819), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(KEYINPUT77), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT2), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n820), .A2(G48), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(G305) );
  NAND2_X1 U681 ( .A1(G49), .A2(n820), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G74), .A2(G651), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n815), .A2(n611), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n612), .A2(G87), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(G288) );
  NAND2_X1 U687 ( .A1(G85), .A2(n816), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G72), .A2(n819), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G60), .A2(n815), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G47), .A2(n820), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(G290) );
  NAND2_X1 U694 ( .A1(G160), .A2(G40), .ZN(n734) );
  INV_X1 U695 ( .A(n734), .ZN(n629) );
  NAND2_X1 U696 ( .A1(G114), .A2(n885), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT84), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G126), .A2(n886), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT83), .B(n622), .Z(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G138), .A2(n881), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G102), .A2(n882), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT64), .ZN(n733) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT91), .Z(n630) );
  INV_X1 U705 ( .A(G1956), .ZN(n937) );
  NOR2_X1 U706 ( .A1(n680), .A2(n937), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n674) );
  NAND2_X1 U708 ( .A1(G65), .A2(n815), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G53), .A2(n820), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G91), .A2(n816), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G78), .A2(n819), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n986) );
  NOR2_X1 U715 ( .A1(n674), .A2(n986), .ZN(n640) );
  INV_X1 U716 ( .A(KEYINPUT28), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n640), .B(n639), .ZN(n678) );
  INV_X1 U718 ( .A(G1996), .ZN(n921) );
  INV_X1 U719 ( .A(KEYINPUT26), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n699), .A2(G1341), .ZN(n663) );
  NAND2_X1 U721 ( .A1(G56), .A2(n815), .ZN(n643) );
  XOR2_X1 U722 ( .A(KEYINPUT14), .B(n643), .Z(n649) );
  NAND2_X1 U723 ( .A1(n816), .A2(G81), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT12), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G68), .A2(n819), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U727 ( .A(KEYINPUT13), .B(n647), .Z(n648) );
  NOR2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n820), .A2(G43), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n992) );
  INV_X1 U731 ( .A(n992), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G54), .A2(n820), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G66), .A2(n815), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G92), .A2(n816), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G79), .A2(n819), .ZN(n656) );
  XNOR2_X1 U737 ( .A(KEYINPUT71), .B(n656), .ZN(n657) );
  NOR2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  OR2_X1 U740 ( .A1(n545), .A2(n992), .ZN(n665) );
  INV_X1 U741 ( .A(n663), .ZN(n664) );
  NOR2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n667), .A2(n666), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n699), .A2(G1348), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(KEYINPUT92), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n680), .A2(G2067), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n986), .A2(n674), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n679), .B(KEYINPUT29), .ZN(n684) );
  XNOR2_X1 U753 ( .A(G1961), .B(KEYINPUT90), .ZN(n957) );
  NAND2_X1 U754 ( .A1(n699), .A2(n957), .ZN(n682) );
  XOR2_X1 U755 ( .A(KEYINPUT25), .B(G2078), .Z(n969) );
  NAND2_X1 U756 ( .A1(n680), .A2(n969), .ZN(n681) );
  NAND2_X1 U757 ( .A1(n682), .A2(n681), .ZN(n690) );
  NOR2_X1 U758 ( .A1(G301), .A2(n690), .ZN(n683) );
  NOR2_X1 U759 ( .A1(n684), .A2(n683), .ZN(n695) );
  NAND2_X1 U760 ( .A1(G8), .A2(n699), .ZN(n698) );
  NOR2_X1 U761 ( .A1(G1966), .A2(n698), .ZN(n706) );
  NOR2_X1 U762 ( .A1(G2084), .A2(n699), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n706), .A2(n707), .ZN(n685) );
  NAND2_X1 U764 ( .A1(G8), .A2(n685), .ZN(n688) );
  INV_X1 U765 ( .A(KEYINPUT30), .ZN(n686) );
  NOR2_X1 U766 ( .A1(n689), .A2(G168), .ZN(n692) );
  AND2_X1 U767 ( .A1(G301), .A2(n690), .ZN(n691) );
  NOR2_X1 U768 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U769 ( .A(n693), .B(KEYINPUT31), .ZN(n694) );
  NOR2_X1 U770 ( .A1(G1971), .A2(n698), .ZN(n701) );
  NOR2_X1 U771 ( .A1(G2090), .A2(n699), .ZN(n700) );
  NOR2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U773 ( .A1(G303), .A2(n702), .ZN(n703) );
  NAND2_X1 U774 ( .A1(G8), .A2(n707), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U776 ( .A(KEYINPUT94), .B(n710), .ZN(n724) );
  NAND2_X1 U777 ( .A1(n725), .A2(n724), .ZN(n714) );
  NAND2_X1 U778 ( .A1(G8), .A2(G166), .ZN(n711) );
  NOR2_X1 U779 ( .A1(G2090), .A2(n711), .ZN(n712) );
  XNOR2_X1 U780 ( .A(n712), .B(KEYINPUT97), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U782 ( .A(n715), .B(KEYINPUT98), .ZN(n716) );
  NOR2_X1 U783 ( .A1(G1981), .A2(G305), .ZN(n717) );
  XOR2_X1 U784 ( .A(n717), .B(KEYINPUT24), .Z(n718) );
  XNOR2_X1 U785 ( .A(KEYINPUT88), .B(n718), .ZN(n719) );
  NOR2_X1 U786 ( .A1(n698), .A2(n719), .ZN(n720) );
  XNOR2_X1 U787 ( .A(KEYINPUT89), .B(n720), .ZN(n721) );
  XOR2_X1 U788 ( .A(G1981), .B(G305), .Z(n998) );
  NAND2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U790 ( .A(n698), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n987), .A2(n722), .ZN(n727) );
  INV_X1 U792 ( .A(n727), .ZN(n723) );
  NOR2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n729) );
  NOR2_X1 U794 ( .A1(G1971), .A2(G303), .ZN(n726) );
  NOR2_X1 U795 ( .A1(n729), .A2(n726), .ZN(n1004) );
  OR2_X1 U796 ( .A1(n727), .A2(n1004), .ZN(n728) );
  NAND2_X1 U797 ( .A1(KEYINPUT33), .A2(n729), .ZN(n730) );
  NOR2_X1 U798 ( .A1(n698), .A2(n730), .ZN(n731) );
  XNOR2_X1 U799 ( .A(n731), .B(KEYINPUT96), .ZN(n732) );
  NOR2_X1 U800 ( .A1(n734), .A2(n733), .ZN(n774) );
  INV_X1 U801 ( .A(n774), .ZN(n761) );
  NAND2_X1 U802 ( .A1(G140), .A2(n881), .ZN(n736) );
  NAND2_X1 U803 ( .A1(G104), .A2(n882), .ZN(n735) );
  NAND2_X1 U804 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U805 ( .A(KEYINPUT34), .B(n737), .ZN(n742) );
  NAND2_X1 U806 ( .A1(G116), .A2(n885), .ZN(n739) );
  NAND2_X1 U807 ( .A1(G128), .A2(n886), .ZN(n738) );
  NAND2_X1 U808 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U809 ( .A(KEYINPUT35), .B(n740), .Z(n741) );
  NOR2_X1 U810 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U811 ( .A(KEYINPUT36), .B(n743), .ZN(n901) );
  XNOR2_X1 U812 ( .A(G2067), .B(KEYINPUT37), .ZN(n772) );
  OR2_X1 U813 ( .A1(n901), .A2(n772), .ZN(n1015) );
  NAND2_X1 U814 ( .A1(G131), .A2(n881), .ZN(n745) );
  NAND2_X1 U815 ( .A1(G107), .A2(n885), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U817 ( .A1(G95), .A2(n882), .ZN(n747) );
  NAND2_X1 U818 ( .A1(G119), .A2(n886), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U821 ( .A(KEYINPUT86), .B(n750), .Z(n895) );
  NAND2_X1 U822 ( .A1(G1991), .A2(n895), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT87), .ZN(n760) );
  NAND2_X1 U824 ( .A1(G141), .A2(n881), .ZN(n753) );
  NAND2_X1 U825 ( .A1(G117), .A2(n885), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n882), .A2(G105), .ZN(n754) );
  XOR2_X1 U828 ( .A(KEYINPUT38), .B(n754), .Z(n755) );
  NOR2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U830 ( .A1(n886), .A2(G129), .ZN(n757) );
  NAND2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n880) );
  AND2_X1 U832 ( .A1(G1996), .A2(n880), .ZN(n759) );
  NOR2_X1 U833 ( .A1(n760), .A2(n759), .ZN(n1027) );
  NOR2_X1 U834 ( .A1(n1027), .A2(n761), .ZN(n768) );
  INV_X1 U835 ( .A(n768), .ZN(n762) );
  XNOR2_X1 U836 ( .A(G1986), .B(G290), .ZN(n994) );
  NOR2_X1 U837 ( .A1(n880), .A2(G1996), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n765), .B(KEYINPUT100), .ZN(n1018) );
  NOR2_X1 U839 ( .A1(G1986), .A2(G290), .ZN(n766) );
  NOR2_X1 U840 ( .A1(G1991), .A2(n895), .ZN(n1024) );
  NOR2_X1 U841 ( .A1(n766), .A2(n1024), .ZN(n767) );
  NOR2_X1 U842 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U843 ( .A1(n1018), .A2(n769), .ZN(n770) );
  XNOR2_X1 U844 ( .A(n770), .B(KEYINPUT39), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n771), .A2(n563), .ZN(n773) );
  NAND2_X1 U846 ( .A1(n901), .A2(n772), .ZN(n1016) );
  NAND2_X1 U847 ( .A1(n773), .A2(n1016), .ZN(n775) );
  NAND2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U849 ( .A(n777), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U850 ( .A(G2443), .B(G2446), .Z(n779) );
  XNOR2_X1 U851 ( .A(G2427), .B(G2451), .ZN(n778) );
  XNOR2_X1 U852 ( .A(n779), .B(n778), .ZN(n785) );
  XOR2_X1 U853 ( .A(G2430), .B(G2454), .Z(n781) );
  XNOR2_X1 U854 ( .A(G1341), .B(G1348), .ZN(n780) );
  XNOR2_X1 U855 ( .A(n781), .B(n780), .ZN(n783) );
  XOR2_X1 U856 ( .A(G2435), .B(G2438), .Z(n782) );
  XNOR2_X1 U857 ( .A(n783), .B(n782), .ZN(n784) );
  XOR2_X1 U858 ( .A(n785), .B(n784), .Z(n786) );
  AND2_X1 U859 ( .A1(G14), .A2(n786), .ZN(G401) );
  NAND2_X1 U860 ( .A1(G135), .A2(n881), .ZN(n788) );
  NAND2_X1 U861 ( .A1(G111), .A2(n885), .ZN(n787) );
  NAND2_X1 U862 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U863 ( .A1(n886), .A2(G123), .ZN(n789) );
  XOR2_X1 U864 ( .A(KEYINPUT18), .B(n789), .Z(n790) );
  NOR2_X1 U865 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U866 ( .A1(n882), .A2(G99), .ZN(n792) );
  NAND2_X1 U867 ( .A1(n793), .A2(n792), .ZN(n1021) );
  XNOR2_X1 U868 ( .A(G2096), .B(n1021), .ZN(n794) );
  OR2_X1 U869 ( .A1(G2100), .A2(n794), .ZN(G156) );
  INV_X1 U870 ( .A(G132), .ZN(G219) );
  INV_X1 U871 ( .A(G82), .ZN(G220) );
  INV_X1 U872 ( .A(G108), .ZN(G238) );
  NAND2_X1 U873 ( .A1(G94), .A2(G452), .ZN(n796) );
  XOR2_X1 U874 ( .A(KEYINPUT68), .B(n796), .Z(G173) );
  NAND2_X1 U875 ( .A1(G7), .A2(G661), .ZN(n797) );
  XNOR2_X1 U876 ( .A(n797), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U877 ( .A(G223), .B(KEYINPUT69), .ZN(n850) );
  NAND2_X1 U878 ( .A1(n850), .A2(G567), .ZN(n798) );
  XOR2_X1 U879 ( .A(KEYINPUT11), .B(n798), .Z(G234) );
  INV_X1 U880 ( .A(G860), .ZN(n806) );
  NOR2_X1 U881 ( .A1(n992), .A2(n806), .ZN(n799) );
  XOR2_X1 U882 ( .A(KEYINPUT70), .B(n799), .Z(G153) );
  NAND2_X1 U883 ( .A1(G868), .A2(G301), .ZN(n801) );
  OR2_X1 U884 ( .A1(n662), .A2(G868), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n801), .A2(n800), .ZN(G284) );
  INV_X1 U886 ( .A(n986), .ZN(G299) );
  NOR2_X1 U887 ( .A1(G868), .A2(G299), .ZN(n804) );
  INV_X1 U888 ( .A(G868), .ZN(n802) );
  NOR2_X1 U889 ( .A1(G286), .A2(n802), .ZN(n803) );
  NOR2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U891 ( .A(KEYINPUT74), .B(n805), .ZN(G297) );
  NAND2_X1 U892 ( .A1(n806), .A2(G559), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n807), .A2(n662), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n808), .B(KEYINPUT75), .ZN(n809) );
  XOR2_X1 U895 ( .A(KEYINPUT16), .B(n809), .Z(G148) );
  NOR2_X1 U896 ( .A1(G868), .A2(n992), .ZN(n812) );
  NAND2_X1 U897 ( .A1(G868), .A2(n662), .ZN(n810) );
  NOR2_X1 U898 ( .A1(G559), .A2(n810), .ZN(n811) );
  NOR2_X1 U899 ( .A1(n812), .A2(n811), .ZN(G282) );
  XNOR2_X1 U900 ( .A(n992), .B(KEYINPUT76), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n662), .A2(G559), .ZN(n813) );
  XNOR2_X1 U902 ( .A(n814), .B(n813), .ZN(n831) );
  NOR2_X1 U903 ( .A1(G860), .A2(n831), .ZN(n825) );
  NAND2_X1 U904 ( .A1(G67), .A2(n815), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G93), .A2(n816), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n824) );
  NAND2_X1 U907 ( .A1(G80), .A2(n819), .ZN(n822) );
  NAND2_X1 U908 ( .A1(G55), .A2(n820), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U910 ( .A1(n824), .A2(n823), .ZN(n834) );
  XNOR2_X1 U911 ( .A(n825), .B(n834), .ZN(G145) );
  XNOR2_X1 U912 ( .A(n986), .B(G288), .ZN(n828) );
  XNOR2_X1 U913 ( .A(G166), .B(n834), .ZN(n826) );
  XNOR2_X1 U914 ( .A(n826), .B(G305), .ZN(n827) );
  XNOR2_X1 U915 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U916 ( .A(KEYINPUT19), .B(n829), .ZN(n830) );
  XNOR2_X1 U917 ( .A(n830), .B(G290), .ZN(n923) );
  XNOR2_X1 U918 ( .A(n831), .B(n923), .ZN(n832) );
  NAND2_X1 U919 ( .A1(n832), .A2(G868), .ZN(n833) );
  XOR2_X1 U920 ( .A(KEYINPUT81), .B(n833), .Z(n836) );
  OR2_X1 U921 ( .A1(n834), .A2(G868), .ZN(n835) );
  NAND2_X1 U922 ( .A1(n836), .A2(n835), .ZN(G295) );
  NAND2_X1 U923 ( .A1(G2078), .A2(G2084), .ZN(n837) );
  XOR2_X1 U924 ( .A(KEYINPUT20), .B(n837), .Z(n838) );
  NAND2_X1 U925 ( .A1(G2090), .A2(n838), .ZN(n839) );
  XNOR2_X1 U926 ( .A(KEYINPUT21), .B(n839), .ZN(n840) );
  NAND2_X1 U927 ( .A1(n840), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U928 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U929 ( .A1(G120), .A2(G69), .ZN(n841) );
  NOR2_X1 U930 ( .A1(G238), .A2(n841), .ZN(n842) );
  NAND2_X1 U931 ( .A1(G57), .A2(n842), .ZN(n856) );
  NAND2_X1 U932 ( .A1(n856), .A2(G567), .ZN(n848) );
  NOR2_X1 U933 ( .A1(G220), .A2(G219), .ZN(n843) );
  XOR2_X1 U934 ( .A(KEYINPUT22), .B(n843), .Z(n844) );
  NOR2_X1 U935 ( .A1(G218), .A2(n844), .ZN(n845) );
  NAND2_X1 U936 ( .A1(G96), .A2(n845), .ZN(n857) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n857), .ZN(n846) );
  XNOR2_X1 U938 ( .A(KEYINPUT82), .B(n846), .ZN(n847) );
  NAND2_X1 U939 ( .A1(n848), .A2(n847), .ZN(n935) );
  NAND2_X1 U940 ( .A1(G483), .A2(G661), .ZN(n849) );
  NOR2_X1 U941 ( .A1(n935), .A2(n849), .ZN(n855) );
  NAND2_X1 U942 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n850), .ZN(G217) );
  NAND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n852) );
  INV_X1 U945 ( .A(G661), .ZN(n851) );
  NOR2_X1 U946 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U947 ( .A(n853), .B(KEYINPUT101), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U949 ( .A1(n855), .A2(n854), .ZN(G188) );
  XOR2_X1 U950 ( .A(G120), .B(KEYINPUT102), .Z(G236) );
  XNOR2_X1 U951 ( .A(G69), .B(KEYINPUT103), .ZN(G235) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  NOR2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n858), .B(KEYINPUT104), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  NAND2_X1 U957 ( .A1(G124), .A2(n886), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G136), .A2(n881), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT106), .B(n860), .Z(n863) );
  NAND2_X1 U961 ( .A1(n882), .A2(G100), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT108), .B(n861), .Z(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G112), .A2(n885), .ZN(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT107), .B(n866), .ZN(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(G162) );
  XNOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n1021), .B(KEYINPUT110), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U971 ( .A(G162), .B(n871), .ZN(n899) );
  NAND2_X1 U972 ( .A1(G118), .A2(n885), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G130), .A2(n886), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n882), .A2(G106), .ZN(n874) );
  XOR2_X1 U976 ( .A(KEYINPUT109), .B(n874), .Z(n876) );
  NAND2_X1 U977 ( .A1(n881), .A2(G142), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n894) );
  XOR2_X1 U981 ( .A(G164), .B(n880), .Z(n892) );
  NAND2_X1 U982 ( .A1(G139), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G103), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n1028) );
  XNOR2_X1 U990 ( .A(n892), .B(n1028), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n897) );
  XNOR2_X1 U992 ( .A(G160), .B(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(n903) );
  XOR2_X1 U997 ( .A(KEYINPUT111), .B(n903), .Z(G395) );
  XOR2_X1 U998 ( .A(G2100), .B(G2096), .Z(n905) );
  XNOR2_X1 U999 ( .A(KEYINPUT42), .B(G2678), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1001 ( .A(KEYINPUT43), .B(G2072), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G2067), .B(G2090), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1005 ( .A(G2078), .B(G2084), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(G227) );
  XOR2_X1 U1007 ( .A(G1956), .B(G1971), .Z(n913) );
  XNOR2_X1 U1008 ( .A(G1991), .B(G1976), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n917) );
  XOR2_X1 U1010 ( .A(G1966), .B(G1961), .Z(n915) );
  XNOR2_X1 U1011 ( .A(G1986), .B(G1981), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n917), .B(n916), .Z(n919) );
  XNOR2_X1 U1014 ( .A(G2474), .B(KEYINPUT105), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(KEYINPUT41), .B(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(G229) );
  XNOR2_X1 U1018 ( .A(n662), .B(n992), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n926) );
  XOR2_X1 U1020 ( .A(G171), .B(G286), .Z(n925) );
  XNOR2_X1 U1021 ( .A(n926), .B(n925), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n927), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(KEYINPUT112), .B(n928), .ZN(G397) );
  NOR2_X1 U1024 ( .A1(G401), .A2(n935), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(G395), .A2(n930), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n933), .A2(G397), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(n934), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(n935), .ZN(G319) );
  INV_X1 U1033 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1034 ( .A(G1348), .B(KEYINPUT59), .Z(n936) );
  XNOR2_X1 U1035 ( .A(G4), .B(n936), .ZN(n944) );
  XOR2_X1 U1036 ( .A(G1981), .B(G6), .Z(n939) );
  XNOR2_X1 U1037 ( .A(n937), .B(G20), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G19), .B(G1341), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(n942), .B(KEYINPUT123), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(KEYINPUT60), .B(n945), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(n946), .B(KEYINPUT124), .ZN(n956) );
  XOR2_X1 U1045 ( .A(G1966), .B(KEYINPUT125), .Z(n947) );
  XNOR2_X1 U1046 ( .A(G21), .B(n947), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G1976), .B(G23), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G1971), .B(G22), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n950) );
  NAND2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G5), .B(n957), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n960), .Z(n961) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n961), .ZN(n1013) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(n962), .B(G34), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(G2084), .B(n963), .ZN(n981) );
  XNOR2_X1 U1062 ( .A(G2090), .B(G35), .ZN(n978) );
  XOR2_X1 U1063 ( .A(G1991), .B(G25), .Z(n964) );
  NAND2_X1 U1064 ( .A1(n964), .A2(G28), .ZN(n975) );
  XOR2_X1 U1065 ( .A(G2072), .B(KEYINPUT117), .Z(n965) );
  XNOR2_X1 U1066 ( .A(G33), .B(n965), .ZN(n967) );
  XNOR2_X1 U1067 ( .A(G26), .B(G2067), .ZN(n966) );
  NOR2_X1 U1068 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1069 ( .A(KEYINPUT118), .B(n968), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G32), .ZN(n971) );
  XNOR2_X1 U1071 ( .A(n969), .B(G27), .ZN(n970) );
  NOR2_X1 U1072 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1075 ( .A(KEYINPUT53), .B(n976), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1077 ( .A(KEYINPUT119), .B(n979), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1079 ( .A(KEYINPUT55), .B(n982), .Z(n983) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n983), .ZN(n1010) );
  XOR2_X1 U1081 ( .A(G16), .B(KEYINPUT56), .Z(n1008) );
  XNOR2_X1 U1082 ( .A(G1348), .B(n662), .ZN(n985) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n984) );
  NAND2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n1006) );
  XNOR2_X1 U1085 ( .A(G1956), .B(n986), .ZN(n988) );
  NAND2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1087 ( .A(G1961), .B(G171), .Z(n989) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n989), .ZN(n990) );
  NOR2_X1 U1089 ( .A1(n991), .A2(n990), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(G168), .B(G1966), .Z(n997) );
  XNOR2_X1 U1094 ( .A(KEYINPUT121), .B(n997), .ZN(n999) );
  NAND2_X1 U1095 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n1000), .Z(n1001) );
  NOR2_X1 U1097 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1011), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT126), .B(n1014), .ZN(n1044) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1038) );
  XOR2_X1 U1106 ( .A(G2090), .B(G162), .Z(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT51), .B(n1019), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(n1020), .B(KEYINPUT115), .ZN(n1036) );
  XNOR2_X1 U1110 ( .A(G160), .B(G2084), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(KEYINPUT114), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1034) );
  XOR2_X1 U1115 ( .A(G2072), .B(n1028), .Z(n1030) );
  XOR2_X1 U1116 ( .A(G164), .B(G2078), .Z(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1118 ( .A(KEYINPUT50), .B(n1031), .Z(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT116), .B(n1032), .ZN(n1033) );
  NOR2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(KEYINPUT52), .B(n1039), .ZN(n1041) );
  INV_X1 U1124 ( .A(KEYINPUT55), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1126 ( .A1(n1042), .A2(G29), .ZN(n1043) );
  NAND2_X1 U1127 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1128 ( .A(n1045), .B(KEYINPUT127), .ZN(n1046) );
  XNOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1046), .ZN(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

