//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND3_X1  g0042(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(new_n216), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G1), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n246), .ZN(new_n251));
  INV_X1    g0051(.A(G107), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT25), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n252), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n250), .A2(G107), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT22), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G87), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT70), .B1(new_n259), .B2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n257), .A2(new_n262), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n248), .A3(KEYINPUT3), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n268), .A2(new_n269), .A3(new_n271), .A4(new_n260), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT23), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT80), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n267), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n272), .A2(new_n273), .B1(new_n277), .B2(G20), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT80), .B1(new_n282), .B2(new_n266), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT24), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n244), .B1(new_n283), .B2(KEYINPUT24), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n256), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n268), .A2(new_n271), .A3(new_n260), .ZN(new_n288));
  INV_X1    g0088(.A(G257), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G250), .B2(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G294), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n291), .B1(new_n248), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT5), .B(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  OAI211_X1 g0097(.A(G1), .B(G13), .C1(new_n248), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n296), .A2(new_n298), .A3(G274), .A4(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n300), .B2(new_n296), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G264), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n295), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G179), .B2(new_n304), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n287), .A2(new_n308), .A3(KEYINPUT81), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT81), .ZN(new_n310));
  INV_X1    g0110(.A(new_n256), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n280), .B1(new_n267), .B2(new_n279), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT24), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n245), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n284), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n310), .B1(new_n315), .B2(new_n307), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(G50), .B1(new_n207), .B2(G1), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n247), .A2(new_n318), .B1(G50), .B2(new_n246), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n207), .A2(G33), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G20), .A2(G33), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n321), .A2(new_n323), .B1(G150), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n203), .A2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n319), .B1(new_n327), .B2(new_n244), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT9), .Z(new_n329));
  INV_X1    g0129(.A(KEYINPUT67), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT3), .B(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G222), .A2(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G223), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n294), .C1(G77), .C2(new_n331), .ZN(new_n336));
  INV_X1    g0136(.A(G226), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n298), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(G1), .B1(new_n297), .B2(new_n299), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n298), .A2(G274), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT65), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n298), .A2(KEYINPUT65), .A3(new_n341), .A4(G274), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n330), .B1(new_n348), .B2(G190), .ZN(new_n349));
  INV_X1    g0149(.A(G200), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n329), .B(new_n349), .C1(new_n350), .C2(new_n348), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT10), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n348), .A2(G169), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n340), .A2(new_n347), .A3(G179), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n353), .A2(new_n328), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n331), .A2(G232), .A3(new_n333), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT66), .B(G107), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(new_n331), .ZN(new_n359));
  INV_X1    g0159(.A(G238), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n261), .A2(new_n360), .A3(new_n333), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n294), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n294), .A2(new_n341), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n344), .A2(new_n345), .B1(G244), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(G179), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G77), .B1(new_n207), .B2(G1), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n247), .A2(new_n368), .B1(G77), .B2(new_n246), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n321), .A2(new_n324), .B1(G20), .B2(G77), .ZN(new_n370));
  XOR2_X1   g0170(.A(KEYINPUT15), .B(G87), .Z(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n372), .B2(new_n322), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n373), .B2(new_n244), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n305), .B2(new_n365), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n374), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(G200), .B2(new_n365), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n352), .A2(new_n356), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n247), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n384));
  INV_X1    g0184(.A(G68), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n324), .A2(G50), .B1(G20), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G77), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n322), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n244), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n251), .A2(new_n385), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT12), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(KEYINPUT11), .A3(new_n244), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n384), .A2(new_n391), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT69), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  MUX2_X1   g0198(.A(G226), .B(G232), .S(G1698), .Z(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n331), .B1(G33), .B2(G97), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n400), .A2(new_n298), .B1(new_n360), .B2(new_n339), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(KEYINPUT68), .B2(new_n346), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT68), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n344), .A2(new_n404), .A3(new_n345), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n346), .A2(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n331), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(new_n294), .B1(G238), .B2(new_n363), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n411), .A3(new_n405), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(G169), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n406), .A2(new_n413), .A3(G179), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n414), .B2(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n398), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n403), .B1(new_n402), .B2(new_n405), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n422));
  OAI21_X1  g0222(.A(G200), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n406), .A2(new_n413), .A3(G190), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n397), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n259), .A2(KEYINPUT70), .A3(G33), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT72), .ZN(new_n431));
  AND2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n268), .A4(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n268), .A2(new_n271), .A3(new_n260), .A4(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT72), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G87), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n333), .A2(G223), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(new_n268), .A3(new_n271), .A4(new_n260), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n433), .A2(new_n435), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n294), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n363), .A2(KEYINPUT74), .A3(G232), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  INV_X1    g0242(.A(G232), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n339), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n441), .A2(new_n444), .B1(new_n344), .B2(new_n345), .ZN(new_n445));
  AOI21_X1  g0245(.A(G200), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT73), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n439), .A2(new_n447), .A3(new_n294), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n439), .B2(new_n294), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n378), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n446), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G58), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n385), .ZN(new_n455));
  OAI21_X1  g0255(.A(G20), .B1(new_n455), .B2(new_n201), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n324), .A2(G159), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT7), .ZN(new_n460));
  AOI21_X1  g0260(.A(G20), .B1(new_n460), .B2(KEYINPUT71), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(KEYINPUT71), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n288), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G68), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n288), .B2(new_n461), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT16), .B(new_n459), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT16), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n460), .B1(new_n331), .B2(G20), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n385), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n458), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n244), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n320), .B1(new_n206), .B2(G20), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n383), .A2(new_n474), .B1(new_n251), .B2(new_n320), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n427), .B1(new_n453), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n440), .A2(KEYINPUT73), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n441), .A2(new_n444), .ZN(new_n479));
  INV_X1    g0279(.A(G179), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(new_n346), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n439), .A2(new_n447), .A3(new_n294), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n440), .A2(new_n445), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n305), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT18), .ZN(new_n487));
  INV_X1    g0287(.A(new_n476), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(KEYINPUT17), .C1(new_n489), .C2(new_n446), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT18), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n483), .A2(new_n476), .A3(new_n491), .A4(new_n485), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n477), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n382), .A2(new_n426), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT4), .A2(G244), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n331), .A2(new_n333), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n268), .A2(new_n271), .A3(G244), .A4(new_n260), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G1698), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT75), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n331), .A2(new_n502), .A3(G250), .A4(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n331), .A2(G250), .A3(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n498), .A2(new_n501), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n294), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n296), .A2(new_n300), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n298), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n301), .B1(new_n509), .B2(new_n289), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n305), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n506), .B2(new_n294), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n480), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n516), .A2(new_n517), .A3(G107), .ZN(new_n518));
  XNOR2_X1  g0318(.A(G97), .B(G107), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n324), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n520), .A2(new_n207), .B1(new_n387), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n358), .B1(new_n469), .B2(new_n470), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n244), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n251), .A2(new_n517), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n250), .A2(G97), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n513), .A2(new_n515), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n514), .A2(G190), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n530), .C1(new_n350), .C2(new_n514), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n358), .A2(new_n262), .A3(new_n517), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n207), .B1(new_n409), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n322), .B2(new_n517), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT78), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n288), .A2(G20), .A3(new_n385), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n244), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n372), .A2(new_n251), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n250), .A2(G87), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n298), .A2(G274), .A3(new_n300), .ZN(new_n546));
  OAI21_X1  g0346(.A(G250), .B1(new_n299), .B2(G1), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n294), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n360), .A2(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n268), .A2(new_n271), .A3(new_n260), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT77), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n500), .A2(new_n333), .B1(new_n248), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n298), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(G200), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT76), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n548), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n551), .B(KEYINPUT77), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n561), .A2(new_n555), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(G190), .C1(new_n562), .C2(new_n298), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n545), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n305), .B1(new_n549), .B2(new_n557), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n560), .B(new_n480), .C1(new_n562), .C2(new_n298), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n250), .A2(new_n371), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n542), .A2(new_n543), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n528), .A2(new_n531), .A3(new_n564), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n304), .A2(new_n350), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G190), .B2(new_n304), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n315), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n289), .A2(new_n333), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G264), .B2(new_n333), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n288), .A2(new_n577), .B1(new_n578), .B2(new_n331), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT79), .ZN(new_n581));
  OAI221_X1 g0381(.A(new_n581), .B1(new_n578), .B2(new_n331), .C1(new_n288), .C2(new_n577), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n298), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n497), .B(new_n207), .C1(G33), .C2(new_n517), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(new_n244), .C1(new_n207), .C2(G116), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n246), .A2(G116), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n250), .B2(G116), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G270), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n301), .B1(new_n509), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n480), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n584), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n583), .A2(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(G169), .A4(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n591), .A2(G169), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n583), .A2(new_n593), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT21), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n595), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n591), .B1(new_n596), .B2(G200), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n378), .B2(new_n596), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n317), .A2(new_n494), .A3(new_n575), .A4(new_n605), .ZN(G372));
  NAND2_X1  g0406(.A1(new_n425), .A2(new_n377), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n420), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n477), .A2(new_n490), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n487), .B(new_n492), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n355), .B1(new_n610), .B2(new_n352), .ZN(new_n611));
  INV_X1    g0411(.A(new_n569), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n564), .A2(new_n569), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n528), .ZN(new_n615));
  INV_X1    g0415(.A(new_n528), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(KEYINPUT26), .A3(new_n569), .A4(new_n564), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n612), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n287), .A2(new_n308), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n602), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n575), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n494), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n611), .A2(new_n623), .ZN(G369));
  NAND3_X1  g0424(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n626), .A2(G213), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G343), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n591), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n605), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n602), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT82), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G330), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n309), .A2(new_n316), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n573), .B1(new_n315), .B2(new_n629), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n619), .B2(new_n629), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n602), .A2(new_n630), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n287), .A2(new_n308), .A3(new_n629), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(G399));
  INV_X1    g0449(.A(new_n210), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G41), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n532), .A2(G116), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G1), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n214), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n602), .A2(new_n309), .A3(new_n316), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n575), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n618), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n657), .B1(new_n660), .B2(new_n629), .ZN(new_n661));
  AOI211_X1 g0461(.A(KEYINPUT29), .B(new_n630), .C1(new_n618), .C2(new_n621), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n512), .A2(new_n480), .A3(new_n304), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n549), .A2(new_n557), .B1(new_n583), .B2(new_n593), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT83), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n549), .A2(new_n557), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n304), .A2(new_n480), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n514), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT83), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n596), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n295), .A2(new_n303), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n514), .A2(new_n584), .A3(new_n675), .A4(new_n594), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n668), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n584), .A2(new_n675), .A3(new_n594), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(KEYINPUT30), .A3(new_n514), .A4(new_n667), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n630), .B1(new_n673), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n677), .B(new_n679), .C1(new_n664), .C2(new_n665), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n629), .A2(new_n682), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n681), .A2(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n575), .A2(new_n605), .A3(new_n317), .A4(new_n629), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n663), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n661), .A2(new_n662), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n656), .B1(new_n688), .B2(G1), .ZN(G364));
  AND2_X1   g0489(.A1(new_n207), .A2(G13), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n206), .B1(new_n690), .B2(G45), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n651), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n210), .A2(new_n331), .ZN(new_n694));
  INV_X1    g0494(.A(G355), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n694), .A2(new_n695), .B1(G116), .B2(new_n210), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n238), .A2(new_n299), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n210), .A2(new_n288), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n299), .B2(new_n215), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n696), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G13), .A2(G33), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT84), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G20), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n216), .B1(G20), .B2(new_n305), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n693), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n207), .A2(new_n480), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G200), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n378), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n378), .A2(G200), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n480), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n710), .A2(G326), .B1(new_n713), .B2(G294), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT87), .Z(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n709), .A2(G190), .ZN(new_n717));
  XNOR2_X1  g0517(.A(KEYINPUT33), .B(G317), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n207), .A2(G179), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n378), .A3(G200), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n717), .A2(new_n718), .B1(new_n721), .B2(G283), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n578), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n708), .A2(new_n711), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT85), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(KEYINPUT85), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(G322), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n719), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n331), .B1(new_n734), .B2(G329), .ZN(new_n735));
  INV_X1    g0535(.A(G311), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n708), .A2(new_n732), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n716), .A2(new_n724), .A3(new_n731), .A4(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT88), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT88), .ZN(new_n741));
  INV_X1    g0541(.A(new_n713), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n517), .ZN(new_n743));
  INV_X1    g0543(.A(new_n717), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(G159), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n385), .B1(new_n745), .B2(KEYINPUT32), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n743), .B(new_n746), .C1(KEYINPUT32), .C2(new_n745), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n331), .B1(new_n723), .B2(new_n262), .C1(new_n252), .C2(new_n720), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT86), .Z(new_n749));
  INV_X1    g0549(.A(new_n710), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n750), .A2(new_n202), .B1(new_n737), .B2(new_n387), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n730), .B2(G58), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n747), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n740), .A2(new_n741), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n707), .B1(new_n754), .B2(new_n704), .ZN(new_n755));
  INV_X1    g0555(.A(new_n703), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n635), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT89), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n637), .A2(new_n693), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n635), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n760), .ZN(G396));
  NAND2_X1  g0561(.A1(new_n622), .A2(new_n629), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n374), .A2(new_n629), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n376), .B1(new_n380), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n377), .A2(new_n629), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT90), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n762), .B(new_n767), .Z(new_n768));
  INV_X1    g0568(.A(new_n687), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n693), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  INV_X1    g0571(.A(new_n704), .ZN(new_n772));
  INV_X1    g0572(.A(new_n701), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n693), .B1(new_n774), .B2(G77), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n744), .A2(new_n776), .B1(new_n723), .B2(new_n252), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G303), .B2(new_n710), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n730), .A2(G294), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n261), .B1(new_n737), .B2(new_n554), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G311), .B2(new_n734), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n743), .B1(G87), .B2(new_n721), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n778), .A2(new_n779), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n721), .A2(G68), .B1(new_n713), .B2(G58), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n202), .B2(new_n723), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n288), .B(new_n785), .C1(G132), .C2(new_n734), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT34), .ZN(new_n787));
  INV_X1    g0587(.A(new_n737), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n710), .A2(G137), .B1(new_n788), .B2(G159), .ZN(new_n789));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  INV_X1    g0590(.A(G143), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n790), .B2(new_n744), .C1(new_n729), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n786), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n783), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n775), .B1(new_n796), .B2(new_n704), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n767), .B2(new_n702), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n771), .A2(new_n798), .ZN(G384));
  INV_X1    g0599(.A(new_n520), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT35), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(KEYINPUT35), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n801), .A2(G116), .A3(new_n217), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT36), .Z(new_n804));
  OR3_X1    g0604(.A1(new_n214), .A2(new_n387), .A3(new_n455), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n202), .A2(G68), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n206), .B(G13), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n467), .A2(new_n244), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n288), .A2(new_n461), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n462), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(G68), .A3(new_n464), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT16), .B1(new_n812), .B2(new_n459), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n475), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(new_n483), .A3(new_n485), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT93), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n453), .C2(new_n476), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n628), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n488), .B1(new_n489), .B2(new_n446), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n816), .B1(new_n820), .B2(new_n815), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT37), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n476), .A2(new_n628), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n820), .A2(new_n823), .A3(new_n486), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n818), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n493), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT92), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n493), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n826), .A2(KEYINPUT38), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT94), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n493), .A2(new_n830), .A3(new_n827), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n830), .B1(new_n493), .B2(new_n827), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n837), .A2(KEYINPUT94), .A3(KEYINPUT38), .A4(new_n826), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n826), .A2(new_n829), .A3(new_n831), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n834), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n820), .A2(new_n486), .A3(new_n824), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT95), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n825), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n825), .A2(new_n845), .ZN(new_n847));
  INV_X1    g0647(.A(new_n493), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n846), .A2(new_n847), .B1(new_n848), .B2(new_n824), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n840), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n832), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT96), .B(KEYINPUT39), .Z(new_n853));
  AOI22_X1  g0653(.A1(new_n842), .A2(KEYINPUT39), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n420), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n629), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n628), .B1(new_n487), .B2(new_n492), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n767), .A2(new_n622), .A3(new_n629), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n765), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n414), .A2(G169), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT14), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n425), .A2(new_n862), .A3(new_n417), .A4(new_n416), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n397), .A2(new_n629), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT91), .ZN(new_n866));
  INV_X1    g0666(.A(new_n864), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n420), .A2(new_n425), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT91), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n863), .A2(new_n869), .A3(new_n864), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n860), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n858), .B1(new_n873), .B2(new_n842), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n857), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n494), .B1(new_n661), .B2(new_n662), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n611), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n875), .B(new_n877), .Z(new_n878));
  NAND2_X1  g0678(.A1(new_n681), .A2(new_n682), .ZN(new_n879));
  OAI211_X1 g0679(.A(KEYINPUT31), .B(new_n630), .C1(new_n673), .C2(new_n680), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n686), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n871), .A2(new_n767), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n851), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT40), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n868), .A2(new_n870), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n869), .B1(new_n863), .B2(new_n864), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n767), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n881), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n842), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n494), .A2(new_n881), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n893), .A2(new_n894), .A3(new_n663), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n878), .A2(new_n895), .B1(new_n206), .B2(new_n690), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n878), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n808), .B1(new_n896), .B2(new_n897), .ZN(G367));
  OR2_X1    g0698(.A1(new_n545), .A2(new_n629), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n569), .A3(new_n564), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n900), .A2(KEYINPUT97), .B1(new_n569), .B2(new_n899), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(KEYINPUT97), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n703), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n705), .B1(new_n210), .B2(new_n372), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n234), .A2(new_n698), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n693), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n750), .A2(new_n791), .B1(new_n723), .B2(new_n454), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n742), .A2(new_n385), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n730), .A2(G150), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n331), .B1(new_n737), .B2(new_n202), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(G137), .B2(new_n734), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n717), .A2(G159), .B1(new_n721), .B2(G77), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n909), .A2(new_n910), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n723), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(G116), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT46), .ZN(new_n917));
  INV_X1    g0717(.A(G317), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n737), .A2(new_n776), .B1(new_n733), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n288), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n917), .B(new_n921), .C1(new_n578), .C2(new_n729), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n710), .A2(G311), .B1(new_n721), .B2(G97), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n923), .B1(new_n292), .B2(new_n744), .C1(new_n358), .C2(new_n742), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n914), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT47), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n906), .B1(new_n926), .B2(new_n704), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n903), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n645), .B1(new_n642), .B2(new_n644), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n636), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n688), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT102), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n929), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n636), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT102), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n688), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n643), .A2(KEYINPUT101), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n616), .A2(new_n630), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n528), .B(new_n531), .C1(new_n530), .C2(new_n629), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n647), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(KEYINPUT99), .B(KEYINPUT44), .Z(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT100), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT100), .ZN(new_n946));
  INV_X1    g0746(.A(new_n940), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n648), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n647), .B2(new_n940), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n943), .A2(new_n946), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n643), .A2(new_n945), .A3(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n932), .A2(new_n936), .A3(new_n937), .A4(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n643), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n945), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT101), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n688), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n651), .B(KEYINPUT41), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n692), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n645), .A2(new_n940), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT42), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n528), .B1(new_n317), .B2(new_n939), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT98), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n629), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n963), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n962), .A2(new_n966), .B1(new_n967), .B2(new_n902), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n902), .A2(new_n967), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n643), .A2(new_n940), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n928), .B1(new_n960), .B2(new_n972), .ZN(G387));
  NAND2_X1  g0773(.A1(new_n934), .A2(new_n688), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n930), .A2(new_n931), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n975), .A3(new_n651), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n642), .A2(new_n756), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n231), .A2(new_n299), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n978), .A2(new_n698), .B1(new_n653), .B2(new_n694), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n320), .A2(KEYINPUT50), .A3(G50), .ZN(new_n980));
  AOI21_X1  g0780(.A(G45), .B1(G68), .B2(G77), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT50), .B1(new_n320), .B2(G50), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n653), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n979), .A2(new_n983), .B1(new_n252), .B2(new_n650), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n693), .B1(new_n984), .B2(new_n706), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n723), .A2(new_n387), .B1(new_n733), .B2(new_n790), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT103), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n920), .B1(new_n517), .B2(new_n720), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT104), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n713), .A2(new_n371), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n385), .B2(new_n737), .ZN(new_n992));
  INV_X1    g0792(.A(G159), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n993), .A2(new_n750), .B1(new_n744), .B2(new_n320), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(G50), .C2(new_n730), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n717), .A2(G311), .B1(new_n788), .B2(G303), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT106), .B(G322), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n750), .B2(new_n998), .C1(new_n729), .C2(new_n918), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n915), .A2(G294), .B1(new_n713), .B2(G283), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT105), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT107), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n920), .B1(G326), .B2(new_n734), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n554), .C2(new_n720), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n996), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n985), .B1(new_n1011), .B2(new_n704), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n934), .A2(new_n692), .B1(new_n977), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n976), .A2(new_n1013), .ZN(G393));
  INV_X1    g0814(.A(new_n956), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n952), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n974), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n651), .C1(new_n953), .C2(new_n957), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT108), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n956), .A2(KEYINPUT108), .A3(new_n952), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n692), .A3(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n705), .B1(new_n517), .B2(new_n210), .C1(new_n241), .C2(new_n698), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n693), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n729), .A2(new_n993), .B1(new_n790), .B2(new_n750), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n742), .A2(new_n387), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n920), .B1(new_n791), .B2(new_n733), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n385), .A2(new_n723), .B1(new_n720), .B2(new_n262), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n717), .A2(G50), .B1(new_n788), .B2(new_n321), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT110), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1027), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n729), .A2(new_n736), .B1(new_n918), .B2(new_n750), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n915), .A2(G283), .B1(new_n713), .B2(G116), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n252), .B2(new_n720), .C1(new_n578), .C2(new_n744), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n261), .B1(new_n737), .B2(new_n292), .C1(new_n733), .C2(new_n998), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1034), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1024), .B1(new_n1042), .B2(new_n704), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n947), .B2(new_n756), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1018), .A2(new_n1022), .A3(new_n1044), .ZN(G390));
  NAND2_X1  g0845(.A1(new_n881), .A2(G330), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n887), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n871), .B1(new_n687), .B2(new_n767), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n860), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n687), .A2(new_n767), .A3(new_n871), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n765), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n630), .B1(new_n618), .B2(new_n659), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n767), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n881), .A2(G330), .A3(new_n767), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1050), .B(new_n1053), .C1(new_n1054), .C2(new_n871), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n494), .A2(new_n881), .A3(G330), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n876), .A2(new_n1057), .A3(new_n611), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n872), .A2(new_n856), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n871), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n851), .A2(new_n856), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n854), .A2(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1047), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n852), .A2(new_n853), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n1069), .A3(new_n1061), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1064), .A2(new_n1063), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n1050), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1060), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1058), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1072), .B(new_n1075), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n651), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G125), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT54), .B(G143), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n331), .B1(new_n733), .B2(new_n1078), .C1(new_n737), .C2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n710), .A2(G128), .B1(new_n713), .B2(G159), .ZN(new_n1081));
  INV_X1    g0881(.A(G137), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1081), .B1(new_n202), .B2(new_n720), .C1(new_n1082), .C2(new_n744), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1080), .B(new_n1083), .C1(G132), .C2(new_n730), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n723), .A2(new_n790), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n744), .A2(new_n358), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1028), .B(new_n1088), .C1(G283), .C2(new_n710), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n261), .B1(new_n733), .B2(new_n292), .C1(new_n517), .C2(new_n737), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n385), .A2(new_n720), .B1(new_n723), .B2(new_n262), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n730), .C2(G116), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1084), .A2(new_n1087), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n693), .B1(new_n321), .B2(new_n774), .C1(new_n1093), .C2(new_n772), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n702), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n854), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n692), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1077), .A2(new_n1098), .ZN(G378));
  OAI21_X1  g0899(.A(new_n693), .B1(new_n774), .B2(G50), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n717), .A2(G132), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1082), .B2(new_n737), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n713), .A2(G150), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n723), .B2(new_n1079), .C1(new_n750), .C2(new_n1078), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(G128), .C2(new_n730), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT59), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n734), .A2(G124), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n248), .A2(new_n297), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT113), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n993), .C2(new_n720), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT114), .Z(new_n1113));
  NAND3_X1  g0913(.A1(new_n1107), .A2(new_n1108), .A3(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n372), .A2(new_n737), .B1(new_n776), .B2(new_n733), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n908), .B(new_n1115), .C1(new_n730), .C2(G107), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n710), .A2(G116), .B1(new_n915), .B2(G77), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n720), .A2(new_n454), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G97), .B2(new_n717), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n920), .A2(G41), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT58), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1120), .A2(G50), .A3(new_n1111), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1114), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1100), .B1(new_n1126), .B2(new_n704), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n352), .A2(new_n356), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n628), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n328), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1128), .B(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1131), .B(new_n1132), .Z(new_n1133));
  OAI21_X1  g0933(.A(new_n1127), .B1(new_n1133), .B2(new_n702), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT115), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1133), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(KEYINPUT40), .A2(new_n883), .B1(new_n842), .B2(new_n889), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n663), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n891), .A2(G330), .A3(new_n1133), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n875), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n857), .A3(new_n1142), .A4(new_n874), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n692), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1076), .A2(new_n1059), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1076), .A2(KEYINPUT117), .A3(new_n1059), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT57), .B1(new_n1153), .B2(new_n1146), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1076), .A2(KEYINPUT117), .A3(new_n1059), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT117), .B1(new_n1076), .B2(new_n1059), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n651), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1148), .B1(new_n1154), .B2(new_n1160), .ZN(G375));
  AOI21_X1  g0961(.A(new_n691), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT118), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1056), .A2(KEYINPUT118), .A3(new_n692), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n693), .B1(new_n774), .B2(G68), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n744), .A2(new_n554), .B1(new_n737), .B2(new_n358), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT119), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n729), .A2(new_n776), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n991), .B1(new_n517), .B2(new_n723), .C1(new_n750), .C2(new_n292), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n261), .B1(new_n733), .B2(new_n578), .C1(new_n387), .C2(new_n720), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1173), .A2(KEYINPUT120), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n744), .A2(new_n1079), .B1(new_n993), .B2(new_n723), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1118), .B(new_n1175), .C1(G132), .C2(new_n710), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n742), .A2(new_n202), .B1(new_n737), .B2(new_n790), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT121), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n730), .A2(G137), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n288), .B1(new_n734), .B2(G128), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1173), .A2(KEYINPUT120), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1174), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1165), .B1(new_n1183), .B2(new_n704), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n871), .B2(new_n773), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1163), .A2(new_n1164), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1049), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1060), .A2(new_n959), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(G381));
  INV_X1    g0989(.A(KEYINPUT122), .ZN(new_n1190));
  INV_X1    g0990(.A(G396), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n976), .A3(new_n1013), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1190), .B1(new_n1194), .B2(G387), .ZN(new_n1195));
  INV_X1    g0995(.A(G378), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n652), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1146), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1155), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1197), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(G387), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1193), .A2(new_n1202), .A3(KEYINPUT122), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1195), .A2(new_n1196), .A3(new_n1201), .A4(new_n1203), .ZN(G407));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1196), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1205), .ZN(G409));
  NAND2_X1  g1006(.A1(G375), .A2(G378), .ZN(new_n1207));
  INV_X1    g1007(.A(G213), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(G343), .ZN(new_n1209));
  AND4_X1   g1009(.A1(new_n1077), .A2(new_n1147), .A3(new_n1098), .A4(new_n1136), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n959), .B(new_n1146), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT126), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1209), .A2(G2897), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1049), .A2(new_n1058), .A3(new_n1055), .A4(KEYINPUT60), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1217), .A2(new_n651), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1187), .B1(new_n1075), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1218), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1186), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1049), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1060), .B2(new_n1219), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1217), .A2(new_n651), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT124), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1218), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(G384), .A3(new_n1186), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1227), .A2(new_n1234), .A3(KEYINPUT125), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1216), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1235), .A2(new_n1216), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1214), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1227), .A2(new_n1234), .A3(KEYINPUT125), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT125), .B1(new_n1227), .B2(new_n1234), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1215), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(KEYINPUT126), .A3(new_n1240), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1213), .A2(new_n1242), .A3(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1018), .A2(new_n1044), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G387), .A2(new_n1022), .A3(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G393), .B(new_n1191), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G390), .B(new_n928), .C1(new_n960), .C2(new_n972), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1252), .A2(new_n1253), .A3(KEYINPUT61), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1212), .B(new_n1255), .C1(new_n1201), .C2(new_n1196), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1209), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1211), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1147), .A2(new_n1077), .A3(new_n1098), .A4(new_n1136), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G375), .B2(G378), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1247), .A2(new_n1254), .A3(new_n1258), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1245), .A2(new_n1240), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1256), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1263), .A2(new_n1255), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1268), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1265), .B1(new_n1274), .B2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(new_n1207), .A2(new_n1205), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1235), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1207), .A2(new_n1205), .A3(new_n1255), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1279), .A2(new_n1275), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1275), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


