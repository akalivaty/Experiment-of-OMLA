//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT81), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT10), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n192), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n196), .A2(KEYINPUT68), .A3(new_n198), .A4(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G143), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n209), .B2(G143), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT69), .B(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n191), .B1(new_n205), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G104), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n217), .A3(G104), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(KEYINPUT84), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G101), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n226), .A2(new_n228), .A3(new_n220), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n229), .A3(KEYINPUT85), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n224), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n228), .A3(new_n220), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n221), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI211_X1 g051(.A(KEYINPUT86), .B(new_n221), .C1(new_n230), .C2(new_n234), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n215), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n196), .A2(new_n240), .A3(new_n198), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n193), .A2(new_n195), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n207), .B1(new_n242), .B2(new_n206), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n241), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n230), .A2(new_n234), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n225), .A2(new_n220), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G101), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT4), .B1(new_n251), .B2(G101), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT65), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G134), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(KEYINPUT65), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(G131), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n258), .A2(new_n262), .A3(new_n267), .A4(new_n263), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n197), .B1(new_n209), .B2(G143), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G128), .B1(new_n207), .B2(new_n211), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n203), .A2(new_n204), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n221), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT85), .B1(new_n225), .B2(new_n229), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n232), .A2(new_n233), .A3(new_n231), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n191), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n239), .A2(new_n255), .A3(new_n270), .A4(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G110), .B(G140), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT82), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n282), .B(new_n284), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n239), .A2(new_n255), .A3(new_n279), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT88), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n269), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n288), .B2(new_n269), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n280), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n278), .A2(KEYINPUT86), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n212), .A2(new_n213), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n296), .A2(new_n210), .B1(new_n203), .B2(new_n204), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n235), .A2(new_n236), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT87), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n274), .A2(new_n278), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n295), .A2(new_n297), .A3(new_n298), .A4(KEYINPUT87), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n269), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT12), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n294), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n285), .B(KEYINPUT83), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(G469), .B(new_n293), .C1(new_n310), .C2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n280), .B1(new_n291), .B2(new_n292), .ZN(new_n319));
  INV_X1    g133(.A(new_n285), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n307), .B(new_n270), .C1(new_n322), .C2(new_n304), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT12), .B1(new_n305), .B2(new_n269), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n287), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI211_X1 g139(.A(G469), .B(G902), .C1(new_n321), .C2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n190), .B1(new_n318), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT97), .B(G475), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G237), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n283), .A3(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n206), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n283), .A3(G143), .A4(G214), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT18), .A2(G131), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G125), .B(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n209), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n338), .B(KEYINPUT80), .Z(new_n339));
  NOR2_X1   g153(.A1(new_n337), .A2(new_n192), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G125), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT78), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n192), .ZN(new_n349));
  OAI211_X1 g163(.A(G146), .B(new_n346), .C1(new_n347), .C2(new_n344), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n334), .B(G131), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(KEYINPUT17), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n334), .A2(KEYINPUT17), .A3(G131), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT96), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n341), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G113), .B(G122), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n219), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n341), .B(new_n357), .C1(new_n352), .C2(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n329), .B1(new_n361), .B2(new_n315), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT19), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n337), .B(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n350), .B1(new_n242), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT95), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n350), .B(new_n367), .C1(new_n242), .C2(new_n364), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n351), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n357), .B1(new_n369), .B2(new_n341), .ZN(new_n370));
  INV_X1    g184(.A(new_n360), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G475), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n376), .B(new_n373), .C1(new_n370), .C2(new_n371), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n362), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n283), .A2(G952), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(G234), .B2(G237), .ZN(new_n380));
  NAND2_X1  g194(.A1(G234), .A2(G237), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(G902), .A3(G953), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT99), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT21), .B(G898), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G478), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n388), .A2(KEYINPUT15), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n206), .A2(G128), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT13), .Z(new_n391));
  NAND2_X1  g205(.A1(new_n213), .A2(G143), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G134), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n256), .A3(new_n390), .ZN(new_n395));
  XOR2_X1   g209(.A(G116), .B(G122), .Z(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G116), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(G122), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n217), .B1(new_n400), .B2(KEYINPUT14), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n401), .A2(new_n396), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n396), .ZN(new_n403));
  INV_X1    g217(.A(new_n395), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n256), .B1(new_n392), .B2(new_n390), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n402), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n398), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n187), .A2(new_n408), .A3(G953), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n406), .A3(new_n409), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n389), .B1(new_n413), .B2(KEYINPUT98), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(KEYINPUT98), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n415), .B2(new_n389), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n378), .A2(new_n387), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G214), .B1(G237), .B2(G902), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n399), .A2(KEYINPUT5), .A3(G119), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n421), .A2(KEYINPUT89), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(KEYINPUT89), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(G113), .A3(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(G116), .B(G119), .Z(new_n425));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT2), .B(G113), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT90), .B(new_n431), .C1(new_n237), .C2(new_n238), .ZN(new_n432));
  INV_X1    g246(.A(new_n430), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n425), .A2(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(KEYINPUT70), .A3(new_n429), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n253), .B2(new_n254), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n295), .A2(new_n298), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT90), .B1(new_n441), .B2(new_n431), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n420), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n431), .B1(new_n237), .B2(new_n238), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(new_n439), .A3(new_n432), .A4(new_n419), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n247), .A2(G125), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT68), .B1(new_n271), .B2(new_n200), .ZN(new_n450));
  INV_X1    g264(.A(new_n204), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n214), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n449), .B1(new_n452), .B2(G125), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n283), .A2(G224), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT92), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n419), .A2(KEYINPUT6), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT91), .B(new_n457), .C1(new_n440), .C2(new_n442), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n446), .A2(new_n439), .A3(new_n432), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT91), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n448), .B(new_n456), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT93), .B(KEYINPUT8), .Z(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n419), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n424), .A2(KEYINPUT94), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n427), .B1(new_n424), .B2(KEYINPUT94), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n430), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n441), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n278), .B1(new_n428), .B2(new_n430), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n454), .A2(KEYINPUT7), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n453), .B(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n474), .B2(new_n447), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n462), .A2(new_n463), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n463), .B1(new_n462), .B2(new_n475), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n417), .B(new_n418), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT100), .B1(new_n327), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n292), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n286), .B1(new_n480), .B2(new_n290), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n280), .B1(new_n323), .B2(new_n324), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n311), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n316), .B1(new_n483), .B2(G469), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n319), .A2(new_n320), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n286), .B1(new_n308), .B2(new_n309), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n314), .B(new_n315), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n189), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT100), .ZN(new_n489));
  INV_X1    g303(.A(new_n418), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n462), .A2(new_n475), .ZN(new_n491));
  INV_X1    g305(.A(new_n463), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n462), .A2(new_n475), .A3(new_n463), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n488), .A2(new_n489), .A3(new_n495), .A4(new_n417), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n338), .B(KEYINPUT80), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n199), .A2(G119), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(G110), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT79), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G110), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n498), .A2(new_n501), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n500), .B1(new_n213), .B2(G119), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT24), .B(G110), .Z(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n350), .B(new_n497), .C1(new_n505), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n349), .A2(new_n350), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n502), .A2(G110), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n315), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n408), .B1(G234), .B2(new_n315), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n520), .A2(new_n521), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n525), .A2(G902), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  INV_X1    g345(.A(G131), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n258), .A2(new_n262), .A3(new_n532), .A4(new_n263), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n260), .A2(new_n263), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(G131), .ZN(new_n536));
  AOI211_X1 g350(.A(KEYINPUT67), .B(new_n532), .C1(new_n260), .C2(new_n263), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n452), .A2(new_n539), .B1(new_n269), .B2(new_n248), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n438), .B1(new_n540), .B2(KEYINPUT30), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n247), .B1(new_n266), .B2(new_n268), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n205), .A2(new_n214), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n533), .B(KEYINPUT71), .C1(new_n536), .C2(new_n537), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT72), .B1(new_n547), .B2(KEYINPUT30), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n544), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n452), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n269), .A2(new_n248), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n550), .A2(KEYINPUT72), .A3(KEYINPUT30), .A4(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n542), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(G101), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G210), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n558), .A2(G237), .A3(G953), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n557), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n564), .A2(KEYINPUT75), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n436), .A2(new_n437), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n550), .A2(new_n551), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n554), .A2(new_n565), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n551), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n541), .B1(new_n572), .B2(new_n552), .ZN(new_n573));
  INV_X1    g387(.A(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n564), .A2(KEYINPUT75), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n569), .B1(new_n576), .B2(new_n566), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n560), .B(new_n561), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT28), .B1(new_n547), .B2(new_n567), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n550), .A2(KEYINPUT28), .A3(new_n551), .A4(new_n567), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n538), .B1(new_n205), .B2(new_n214), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n438), .B1(new_n582), .B2(new_n543), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT28), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n568), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n583), .A3(new_n581), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n578), .B1(new_n589), .B2(new_n579), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n531), .B1(new_n577), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT32), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n554), .A2(new_n568), .A3(new_n565), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT31), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n579), .B1(new_n580), .B2(new_n584), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n585), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n598), .A3(new_n569), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT32), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n531), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n573), .A2(new_n574), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n579), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n589), .A2(new_n564), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT29), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n550), .A2(new_n551), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n438), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT77), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n568), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(KEYINPUT77), .A3(new_n438), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT28), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n588), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n564), .A2(KEYINPUT29), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n315), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n606), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n530), .B1(new_n602), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n479), .A2(new_n496), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n226), .A2(new_n228), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G3));
  INV_X1    g434(.A(new_n530), .ZN(new_n621));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n599), .B2(new_n315), .ZN(new_n623));
  INV_X1    g437(.A(new_n531), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n575), .A2(KEYINPUT31), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n594), .A2(KEYINPUT31), .B1(new_n603), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n626), .B2(new_n598), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n488), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n418), .B(new_n387), .C1(new_n476), .C2(new_n477), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n411), .A2(new_n412), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n411), .A2(KEYINPUT101), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n411), .B(new_n412), .C1(KEYINPUT101), .C2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(G478), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n388), .A2(new_n315), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n413), .B2(new_n388), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n378), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT102), .B1(new_n631), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n495), .A2(new_n641), .A3(new_n644), .A4(new_n387), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n630), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n375), .A2(new_n377), .ZN(new_n649));
  INV_X1    g463(.A(new_n362), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n631), .A2(new_n651), .A3(new_n416), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n630), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G107), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT103), .B(KEYINPUT35), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n515), .B(new_n657), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n524), .A2(new_n525), .B1(new_n528), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n623), .A2(new_n627), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n479), .A2(new_n496), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AOI21_X1  g477(.A(new_n659), .B1(new_n602), .B2(new_n616), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n383), .A2(G900), .ZN(new_n665));
  INV_X1    g479(.A(new_n380), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n651), .A2(new_n416), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n495), .A2(KEYINPUT104), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n418), .B1(new_n476), .B2(new_n477), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n651), .A2(new_n416), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n667), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n664), .A2(new_n488), .A3(new_n670), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n667), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n488), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT40), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n493), .A2(new_n494), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT38), .Z(new_n682));
  AND2_X1   g496(.A1(new_n610), .A2(new_n611), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n315), .B1(new_n683), .B2(new_n564), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n603), .A2(new_n579), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(KEYINPUT32), .B(new_n624), .C1(new_n626), .C2(new_n598), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n600), .B1(new_n599), .B2(new_n531), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n659), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n378), .A2(new_n416), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n418), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n682), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n680), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT105), .B(G143), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G45));
  NOR3_X1   g510(.A1(new_n378), .A2(new_n640), .A3(new_n668), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n418), .C1(new_n476), .C2(new_n477), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n616), .B1(new_n687), .B2(new_n688), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n658), .A2(new_n528), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n526), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n699), .A2(new_n700), .A3(new_n488), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NAND2_X1  g518(.A1(new_n308), .A2(new_n309), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n705), .A2(new_n287), .B1(new_n319), .B2(new_n320), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n487), .A3(new_n190), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n617), .A2(new_n643), .A3(new_n645), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND3_X1  g526(.A1(new_n617), .A2(new_n652), .A3(new_n709), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  INV_X1    g528(.A(new_n478), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n664), .A2(new_n715), .A3(new_n709), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  OAI211_X1 g531(.A(new_n418), .B(new_n691), .C1(new_n476), .C2(new_n477), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n613), .A2(new_n579), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n624), .B1(new_n626), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n623), .A2(new_n530), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n709), .A2(new_n719), .A3(new_n387), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NOR2_X1   g538(.A1(new_n708), .A2(new_n672), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n315), .B1(new_n577), .B2(new_n591), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n720), .A2(new_n595), .A3(new_n569), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n726), .A2(G472), .B1(new_n531), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n728), .B2(new_n702), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n623), .A2(new_n721), .A3(new_n659), .A4(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n725), .B(new_n697), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NOR4_X1   g547(.A1(new_n476), .A2(new_n477), .A3(new_n189), .A4(new_n490), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n318), .B2(new_n326), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n484), .A2(KEYINPUT107), .A3(new_n487), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(KEYINPUT42), .A3(new_n617), .A4(new_n697), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n700), .A2(new_n621), .A3(new_n697), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  AND2_X1   g559(.A1(new_n736), .A2(new_n737), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n617), .A3(new_n669), .A4(new_n734), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  AND2_X1   g562(.A1(new_n483), .A2(KEYINPUT45), .ZN(new_n749));
  OAI21_X1  g563(.A(G469), .B1(new_n483), .B2(KEYINPUT45), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n317), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n326), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n752), .B2(new_n751), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n190), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n678), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n651), .A2(KEYINPUT43), .A3(new_n640), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT43), .B1(new_n651), .B2(new_n640), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n702), .A3(new_n758), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(new_n628), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n681), .A2(new_n490), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n756), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  NAND2_X1  g582(.A1(new_n755), .A2(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n754), .A2(new_n190), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n697), .ZN(new_n774));
  OR4_X1    g588(.A1(new_n700), .A2(new_n765), .A3(new_n621), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n342), .ZN(G42));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n707), .A2(new_n487), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n773), .B1(new_n190), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n757), .A2(new_n380), .A3(new_n758), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n722), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n764), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n784), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n682), .A2(new_n490), .A3(new_n709), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n765), .A2(new_n708), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT115), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n783), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n729), .B2(new_n731), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n530), .A2(new_n666), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n792), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n689), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n378), .A3(new_n640), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n789), .A2(new_n790), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n791), .A2(new_n798), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n778), .B1(new_n786), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n804), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n379), .B1(new_n784), .B2(new_n725), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n800), .A2(new_n641), .A3(new_n801), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n797), .B2(new_n617), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n617), .ZN(new_n816));
  AOI211_X1 g630(.A(KEYINPUT117), .B(new_n816), .C1(new_n794), .C2(new_n796), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n818), .A3(KEYINPUT48), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT48), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n814), .B2(new_n817), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n812), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT118), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(KEYINPUT118), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n805), .B(new_n807), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n739), .A2(new_n743), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n710), .A2(new_n713), .A3(new_n716), .A4(new_n723), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n564), .B1(new_n612), .B2(new_n588), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n531), .B1(new_n577), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(G902), .B1(new_n626), .B2(new_n598), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n702), .B(new_n829), .C1(new_n830), .C2(new_n622), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n730), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n726), .A2(G472), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(KEYINPUT106), .A3(new_n702), .A4(new_n829), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n774), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n738), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n378), .A2(new_n416), .A3(new_n667), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n664), .A2(new_n488), .A3(new_n764), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n747), .A3(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n826), .A2(new_n827), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n631), .A2(new_n642), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n628), .A3(new_n621), .A4(new_n488), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n618), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n618), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n653), .A2(new_n661), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n675), .A2(new_n670), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n700), .A2(new_n488), .A3(new_n702), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n848), .A2(new_n849), .B1(new_n835), .B2(new_n725), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n668), .A2(new_n189), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n719), .A2(new_n736), .A3(new_n737), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n703), .B1(new_n852), .B2(new_n690), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n854), .A3(KEYINPUT52), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n676), .A2(new_n732), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n856), .B1(new_n857), .B2(new_n853), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n840), .A2(new_n847), .A3(new_n859), .A4(KEYINPUT53), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n836), .A2(new_n747), .A3(new_n838), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n710), .A2(new_n713), .A3(new_n716), .A4(new_n723), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n744), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n618), .A2(new_n843), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT108), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n618), .A2(new_n841), .A3(new_n843), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n653), .A2(new_n661), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(KEYINPUT111), .A3(KEYINPUT53), .A4(new_n859), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n855), .A2(KEYINPUT109), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT109), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n850), .A2(new_n854), .A3(new_n875), .A4(KEYINPUT52), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n702), .B1(new_n602), .B2(new_n686), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n746), .A2(new_n877), .A3(new_n719), .A4(new_n851), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n676), .A3(new_n732), .A4(new_n703), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n856), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n879), .B2(new_n856), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n874), .B(new_n876), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n883), .B2(new_n871), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n864), .A2(KEYINPUT112), .A3(new_n744), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT112), .B1(new_n864), .B2(new_n744), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n870), .A2(new_n889), .A3(new_n839), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n840), .A2(new_n847), .A3(new_n859), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n889), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n825), .A2(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n651), .A2(new_n640), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n621), .A2(new_n190), .A3(new_n418), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n779), .B2(KEYINPUT49), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n682), .A2(new_n900), .A3(new_n801), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(G75));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n891), .A2(new_n893), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G902), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n558), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n448), .B1(new_n459), .B2(new_n461), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n456), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT55), .Z(new_n910));
  AND2_X1   g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n907), .A2(new_n910), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n283), .A2(G952), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G51));
  NAND2_X1  g728(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n895), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n316), .B(KEYINPUT57), .Z(new_n918));
  OAI22_X1  g732(.A1(new_n917), .A2(new_n918), .B1(new_n485), .B2(new_n486), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n906), .A2(new_n749), .A3(new_n750), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n913), .B1(new_n919), .B2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT119), .Z(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n905), .A2(G902), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n913), .B1(new_n925), .B2(new_n372), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n372), .B2(new_n925), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n926), .B(KEYINPUT120), .C1(new_n372), .C2(new_n925), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(G60));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n634), .A2(new_n636), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n638), .B(KEYINPUT59), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n896), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n933), .A2(new_n935), .ZN(new_n938));
  INV_X1    g752(.A(new_n895), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n894), .B1(new_n891), .B2(new_n893), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n913), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n932), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n913), .B1(new_n916), .B2(new_n938), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n885), .B2(new_n895), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n945), .B(KEYINPUT121), .C1(new_n934), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT122), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT60), .Z(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n891), .B2(new_n893), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n913), .B1(new_n952), .B2(new_n658), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n527), .B(KEYINPUT123), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G66));
  INV_X1    g772(.A(new_n385), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n283), .B1(new_n959), .B2(G224), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n870), .A2(new_n827), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n962), .B2(new_n283), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n908), .B1(G898), .B2(new_n283), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(G69));
  AOI21_X1  g779(.A(new_n857), .B1(new_n849), .B2(new_n699), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n767), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n767), .A2(new_n969), .A3(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n756), .A2(new_n617), .A3(new_n719), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n744), .A3(new_n747), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n776), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n974), .A3(new_n283), .ZN(new_n975));
  OAI22_X1  g789(.A1(new_n548), .A2(new_n553), .B1(KEYINPUT30), .B2(new_n540), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(new_n364), .Z(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(G900), .B2(G953), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n773), .A2(new_n775), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n966), .A2(new_n694), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n764), .B1(new_n641), .B2(new_n673), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n816), .A2(new_n983), .A3(new_n679), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n756), .B2(new_n766), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n283), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n977), .B(KEYINPUT124), .Z(new_n988));
  AOI22_X1  g802(.A1(new_n975), .A2(new_n978), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(G72));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n986), .B2(new_n962), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n913), .B1(new_n994), .B2(new_n685), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n971), .A2(new_n974), .A3(new_n961), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n993), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n604), .B(KEYINPUT126), .Z(new_n998));
  OAI21_X1  g812(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n604), .A2(new_n993), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n685), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n873), .B2(new_n884), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n999), .B1(new_n1003), .B2(new_n1004), .ZN(G57));
endmodule


