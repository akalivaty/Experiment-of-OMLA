

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U545 ( .A(n682), .B(n681), .ZN(n761) );
  AND2_X1 U546 ( .A1(n800), .A2(n747), .ZN(n751) );
  AND2_X1 U547 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X2 U548 ( .A1(n684), .A2(n762), .ZN(n729) );
  NOR2_X1 U549 ( .A1(n723), .A2(n722), .ZN(n725) );
  XNOR2_X1 U550 ( .A(KEYINPUT99), .B(n717), .ZN(n745) );
  XNOR2_X1 U551 ( .A(n761), .B(n683), .ZN(n684) );
  INV_X1 U552 ( .A(KEYINPUT96), .ZN(n683) );
  XNOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT32), .ZN(n738) );
  INV_X1 U554 ( .A(KEYINPUT64), .ZN(n753) );
  INV_X1 U555 ( .A(KEYINPUT27), .ZN(n690) );
  XNOR2_X1 U556 ( .A(n691), .B(n690), .ZN(n693) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n695) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n724) );
  XNOR2_X1 U559 ( .A(n739), .B(n738), .ZN(n800) );
  NAND2_X1 U560 ( .A1(G8), .A2(n729), .ZN(n807) );
  INV_X1 U561 ( .A(KEYINPUT105), .ZN(n815) );
  INV_X1 U562 ( .A(G2104), .ZN(n532) );
  NOR2_X2 U563 ( .A1(n536), .A2(n532), .ZN(n894) );
  NOR2_X1 U564 ( .A1(G651), .A2(n638), .ZN(n646) );
  NOR2_X1 U565 ( .A1(n541), .A2(n540), .ZN(n680) );
  XOR2_X1 U566 ( .A(G2443), .B(G2446), .Z(n513) );
  XNOR2_X1 U567 ( .A(G2427), .B(G2451), .ZN(n512) );
  XNOR2_X1 U568 ( .A(n513), .B(n512), .ZN(n519) );
  XOR2_X1 U569 ( .A(G2430), .B(G2454), .Z(n515) );
  XNOR2_X1 U570 ( .A(G1341), .B(G1348), .ZN(n514) );
  XNOR2_X1 U571 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U572 ( .A(G2435), .B(G2438), .Z(n516) );
  XNOR2_X1 U573 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U574 ( .A(n519), .B(n518), .Z(n520) );
  AND2_X1 U575 ( .A1(G14), .A2(n520), .ZN(G401) );
  INV_X1 U576 ( .A(G651), .ZN(n525) );
  NOR2_X1 U577 ( .A1(G543), .A2(n525), .ZN(n521) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n521), .Z(n645) );
  NAND2_X1 U579 ( .A1(G64), .A2(n645), .ZN(n523) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n638) );
  NAND2_X1 U581 ( .A1(G52), .A2(n646), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U583 ( .A(KEYINPUT69), .B(n524), .Z(n531) );
  OR2_X1 U584 ( .A1(n525), .A2(n638), .ZN(n526) );
  XNOR2_X1 U585 ( .A(KEYINPUT65), .B(n526), .ZN(n641) );
  NAND2_X1 U586 ( .A1(G77), .A2(n641), .ZN(n528) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U588 ( .A1(G90), .A2(n642), .ZN(n527) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U590 ( .A(KEYINPUT9), .B(n529), .Z(n530) );
  NOR2_X1 U591 ( .A1(n531), .A2(n530), .ZN(G171) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G69), .ZN(G235) );
  INV_X1 U594 ( .A(G108), .ZN(G238) );
  INV_X1 U595 ( .A(G120), .ZN(G236) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  INV_X1 U598 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n894), .A2(G113), .ZN(n535) );
  NOR2_X1 U600 ( .A1(G2105), .A2(n532), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G101), .A2(n542), .ZN(n533) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U603 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X2 U604 ( .A1(G2104), .A2(n536), .ZN(n895) );
  NAND2_X1 U605 ( .A1(G125), .A2(n895), .ZN(n539) );
  NOR2_X1 U606 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X1 U607 ( .A(KEYINPUT17), .B(n537), .Z(n601) );
  NAND2_X1 U608 ( .A1(G137), .A2(n601), .ZN(n538) );
  NAND2_X1 U609 ( .A1(n539), .A2(n538), .ZN(n540) );
  BUF_X1 U610 ( .A(n680), .Z(G160) );
  BUF_X1 U611 ( .A(n542), .Z(n898) );
  NAND2_X1 U612 ( .A1(G102), .A2(n898), .ZN(n544) );
  NAND2_X1 U613 ( .A1(G138), .A2(n601), .ZN(n543) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G114), .A2(n894), .ZN(n546) );
  NAND2_X1 U616 ( .A1(G126), .A2(n895), .ZN(n545) );
  NAND2_X1 U617 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U618 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U619 ( .A1(G63), .A2(n645), .ZN(n550) );
  NAND2_X1 U620 ( .A1(G51), .A2(n646), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(n551), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n642), .A2(G89), .ZN(n552) );
  XNOR2_X1 U624 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U625 ( .A1(G76), .A2(n641), .ZN(n553) );
  NAND2_X1 U626 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U627 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  NOR2_X1 U628 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U629 ( .A(KEYINPUT75), .B(n558), .Z(n559) );
  XOR2_X1 U630 ( .A(KEYINPUT7), .B(n559), .Z(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n560) );
  XOR2_X1 U633 ( .A(n560), .B(KEYINPUT10), .Z(n917) );
  NAND2_X1 U634 ( .A1(n917), .A2(G567), .ZN(n561) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n561), .Z(G234) );
  XOR2_X1 U636 ( .A(G860), .B(KEYINPUT74), .Z(n592) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n563) );
  NAND2_X1 U638 ( .A1(G56), .A2(n645), .ZN(n562) );
  XNOR2_X1 U639 ( .A(n563), .B(n562), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G81), .A2(n642), .ZN(n564) );
  XOR2_X1 U641 ( .A(KEYINPUT12), .B(n564), .Z(n565) );
  XNOR2_X1 U642 ( .A(n565), .B(KEYINPUT73), .ZN(n567) );
  NAND2_X1 U643 ( .A1(G68), .A2(n641), .ZN(n566) );
  NAND2_X1 U644 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n568), .Z(n569) );
  NOR2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n646), .A2(G43), .ZN(n571) );
  NAND2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n938) );
  OR2_X1 U649 ( .A1(n592), .A2(n938), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G79), .A2(n641), .ZN(n574) );
  NAND2_X1 U653 ( .A1(G54), .A2(n646), .ZN(n573) );
  NAND2_X1 U654 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U655 ( .A1(G92), .A2(n642), .ZN(n576) );
  NAND2_X1 U656 ( .A1(G66), .A2(n645), .ZN(n575) );
  NAND2_X1 U657 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U659 ( .A(n579), .B(KEYINPUT15), .Z(n925) );
  INV_X1 U660 ( .A(n925), .ZN(n839) );
  INV_X1 U661 ( .A(G868), .ZN(n662) );
  NAND2_X1 U662 ( .A1(n839), .A2(n662), .ZN(n580) );
  NAND2_X1 U663 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n642), .ZN(n583) );
  NAND2_X1 U665 ( .A1(G65), .A2(n645), .ZN(n582) );
  NAND2_X1 U666 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n646), .A2(G53), .ZN(n584) );
  XOR2_X1 U668 ( .A(KEYINPUT70), .B(n584), .Z(n585) );
  NOR2_X1 U669 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n641), .A2(G78), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n588), .A2(n587), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n662), .ZN(n589) );
  XNOR2_X1 U673 ( .A(n589), .B(KEYINPUT76), .ZN(n591) );
  NOR2_X1 U674 ( .A1(G299), .A2(G868), .ZN(n590) );
  NOR2_X1 U675 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n592), .A2(G559), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n593), .A2(n925), .ZN(n594) );
  XNOR2_X1 U678 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n938), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n925), .A2(G868), .ZN(n595) );
  NOR2_X1 U681 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U682 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G99), .A2(n898), .ZN(n599) );
  NAND2_X1 U684 ( .A1(G111), .A2(n894), .ZN(n598) );
  NAND2_X1 U685 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U686 ( .A(n600), .B(KEYINPUT77), .ZN(n603) );
  BUF_X1 U687 ( .A(n601), .Z(n900) );
  NAND2_X1 U688 ( .A1(G135), .A2(n900), .ZN(n602) );
  NAND2_X1 U689 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n895), .A2(G123), .ZN(n604) );
  XOR2_X1 U691 ( .A(KEYINPUT18), .B(n604), .Z(n605) );
  NOR2_X1 U692 ( .A1(n606), .A2(n605), .ZN(n990) );
  XOR2_X1 U693 ( .A(G2096), .B(n990), .Z(n607) );
  NOR2_X1 U694 ( .A1(G2100), .A2(n607), .ZN(n608) );
  XOR2_X1 U695 ( .A(KEYINPUT78), .B(n608), .Z(G156) );
  NAND2_X1 U696 ( .A1(G93), .A2(n642), .ZN(n610) );
  NAND2_X1 U697 ( .A1(G67), .A2(n645), .ZN(n609) );
  NAND2_X1 U698 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U699 ( .A1(G80), .A2(n641), .ZN(n612) );
  NAND2_X1 U700 ( .A1(G55), .A2(n646), .ZN(n611) );
  NAND2_X1 U701 ( .A1(n612), .A2(n611), .ZN(n613) );
  OR2_X1 U702 ( .A1(n614), .A2(n613), .ZN(n661) );
  NAND2_X1 U703 ( .A1(G559), .A2(n925), .ZN(n615) );
  XNOR2_X1 U704 ( .A(n615), .B(n938), .ZN(n658) );
  NOR2_X1 U705 ( .A1(G860), .A2(n658), .ZN(n616) );
  XOR2_X1 U706 ( .A(KEYINPUT79), .B(n616), .Z(n617) );
  XOR2_X1 U707 ( .A(n661), .B(n617), .Z(G145) );
  NAND2_X1 U708 ( .A1(G86), .A2(n642), .ZN(n619) );
  NAND2_X1 U709 ( .A1(G61), .A2(n645), .ZN(n618) );
  NAND2_X1 U710 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U711 ( .A(KEYINPUT80), .B(n620), .ZN(n623) );
  NAND2_X1 U712 ( .A1(n641), .A2(G73), .ZN(n621) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n621), .Z(n622) );
  NOR2_X1 U714 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n646), .A2(G48), .ZN(n624) );
  NAND2_X1 U716 ( .A1(n625), .A2(n624), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G60), .A2(n645), .ZN(n627) );
  NAND2_X1 U718 ( .A1(G47), .A2(n646), .ZN(n626) );
  NAND2_X1 U719 ( .A1(n627), .A2(n626), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n641), .A2(G72), .ZN(n628) );
  XNOR2_X1 U721 ( .A(n628), .B(KEYINPUT66), .ZN(n630) );
  NAND2_X1 U722 ( .A1(G85), .A2(n642), .ZN(n629) );
  NAND2_X1 U723 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U724 ( .A(KEYINPUT67), .B(n631), .Z(n632) );
  NOR2_X1 U725 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U726 ( .A(KEYINPUT68), .B(n634), .Z(G290) );
  NAND2_X1 U727 ( .A1(G49), .A2(n646), .ZN(n636) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U729 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U730 ( .A1(n645), .A2(n637), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U732 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U733 ( .A1(G75), .A2(n641), .ZN(n644) );
  NAND2_X1 U734 ( .A1(G88), .A2(n642), .ZN(n643) );
  NAND2_X1 U735 ( .A1(n644), .A2(n643), .ZN(n650) );
  NAND2_X1 U736 ( .A1(G62), .A2(n645), .ZN(n648) );
  NAND2_X1 U737 ( .A1(G50), .A2(n646), .ZN(n647) );
  NAND2_X1 U738 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U739 ( .A1(n650), .A2(n649), .ZN(G166) );
  INV_X1 U740 ( .A(G166), .ZN(G303) );
  XOR2_X1 U741 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n652) );
  XOR2_X1 U742 ( .A(G299), .B(KEYINPUT82), .Z(n651) );
  XNOR2_X1 U743 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U744 ( .A(n661), .B(n653), .Z(n655) );
  XOR2_X1 U745 ( .A(G288), .B(G303), .Z(n654) );
  XNOR2_X1 U746 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U747 ( .A(G290), .B(n656), .Z(n657) );
  XNOR2_X1 U748 ( .A(G305), .B(n657), .ZN(n840) );
  XNOR2_X1 U749 ( .A(KEYINPUT83), .B(n658), .ZN(n659) );
  XNOR2_X1 U750 ( .A(n840), .B(n659), .ZN(n660) );
  NAND2_X1 U751 ( .A1(n660), .A2(G868), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U753 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U760 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U763 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U764 ( .A1(G96), .A2(n671), .ZN(n837) );
  NAND2_X1 U765 ( .A1(n837), .A2(G2106), .ZN(n676) );
  NOR2_X1 U766 ( .A1(G237), .A2(G236), .ZN(n673) );
  NOR2_X1 U767 ( .A1(G238), .A2(G235), .ZN(n672) );
  NAND2_X1 U768 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U769 ( .A(KEYINPUT84), .B(n674), .ZN(n838) );
  NAND2_X1 U770 ( .A1(n838), .A2(G567), .ZN(n675) );
  NAND2_X1 U771 ( .A1(n676), .A2(n675), .ZN(n916) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n677) );
  XOR2_X1 U773 ( .A(KEYINPUT85), .B(n677), .Z(n678) );
  NOR2_X1 U774 ( .A1(n916), .A2(n678), .ZN(n836) );
  NAND2_X1 U775 ( .A1(n836), .A2(G36), .ZN(n679) );
  XNOR2_X1 U776 ( .A(KEYINPUT86), .B(n679), .ZN(G176) );
  NAND2_X1 U777 ( .A1(n680), .A2(G40), .ZN(n682) );
  INV_X1 U778 ( .A(KEYINPUT87), .ZN(n681) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n762) );
  XOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .Z(n971) );
  NOR2_X1 U781 ( .A1(n971), .A2(n729), .ZN(n685) );
  XOR2_X1 U782 ( .A(KEYINPUT100), .B(n685), .Z(n687) );
  INV_X1 U783 ( .A(G1961), .ZN(n860) );
  NAND2_X1 U784 ( .A1(n729), .A2(n860), .ZN(n686) );
  NAND2_X1 U785 ( .A1(n687), .A2(n686), .ZN(n721) );
  AND2_X1 U786 ( .A1(n721), .A2(G171), .ZN(n688) );
  XNOR2_X1 U787 ( .A(n688), .B(KEYINPUT101), .ZN(n716) );
  INV_X1 U788 ( .A(G299), .ZN(n698) );
  INV_X1 U789 ( .A(n729), .ZN(n689) );
  NAND2_X1 U790 ( .A1(n689), .A2(G2072), .ZN(n691) );
  NAND2_X1 U791 ( .A1(G1956), .A2(n729), .ZN(n692) );
  NAND2_X1 U792 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U793 ( .A(n694), .B(KEYINPUT102), .Z(n697) );
  NOR2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n696) );
  XNOR2_X1 U795 ( .A(n696), .B(n695), .ZN(n713) );
  NAND2_X1 U796 ( .A1(n698), .A2(n697), .ZN(n711) );
  AND2_X1 U797 ( .A1(n689), .A2(G1996), .ZN(n699) );
  XOR2_X1 U798 ( .A(n699), .B(KEYINPUT26), .Z(n701) );
  NAND2_X1 U799 ( .A1(n729), .A2(G1341), .ZN(n700) );
  NAND2_X1 U800 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U801 ( .A1(n938), .A2(n702), .ZN(n706) );
  NAND2_X1 U802 ( .A1(G1348), .A2(n729), .ZN(n704) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n689), .ZN(n703) );
  NAND2_X1 U804 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U805 ( .A1(n839), .A2(n707), .ZN(n705) );
  OR2_X1 U806 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n839), .A2(n707), .ZN(n708) );
  NAND2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U811 ( .A(n714), .B(KEYINPUT29), .Z(n715) );
  NAND2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n729), .ZN(n741) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n807), .ZN(n717) );
  NAND2_X1 U815 ( .A1(G8), .A2(n745), .ZN(n718) );
  NOR2_X1 U816 ( .A1(n741), .A2(n718), .ZN(n719) );
  XOR2_X1 U817 ( .A(KEYINPUT30), .B(n719), .Z(n720) );
  NOR2_X1 U818 ( .A1(G168), .A2(n720), .ZN(n723) );
  NOR2_X1 U819 ( .A1(G171), .A2(n721), .ZN(n722) );
  XNOR2_X1 U820 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n740) );
  AND2_X1 U822 ( .A1(G286), .A2(G8), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n740), .A2(n728), .ZN(n737) );
  INV_X1 U824 ( .A(G8), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n807), .ZN(n731) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U828 ( .A(KEYINPUT103), .B(n732), .Z(n733) );
  NAND2_X1 U829 ( .A1(n733), .A2(G303), .ZN(n734) );
  OR2_X1 U830 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U831 ( .A(n740), .ZN(n744) );
  NAND2_X1 U832 ( .A1(G8), .A2(n741), .ZN(n742) );
  XOR2_X1 U833 ( .A(KEYINPUT98), .B(n742), .Z(n743) );
  NOR2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n799) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n921) );
  AND2_X1 U837 ( .A1(n799), .A2(n921), .ZN(n747) );
  INV_X1 U838 ( .A(n921), .ZN(n749) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n757), .A2(n748), .ZN(n922) );
  NOR2_X1 U842 ( .A1(n749), .A2(n922), .ZN(n750) );
  NOR2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n807), .A2(n752), .ZN(n754) );
  XNOR2_X1 U845 ( .A(n754), .B(n753), .ZN(n756) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n755) );
  AND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U849 ( .A1(n758), .A2(n807), .ZN(n759) );
  NOR2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n798) );
  XOR2_X1 U851 ( .A(G1981), .B(G305), .Z(n933) );
  NOR2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n829) );
  XOR2_X1 U853 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n776) );
  NAND2_X1 U854 ( .A1(n900), .A2(G140), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n763), .B(KEYINPUT88), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G104), .A2(n898), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n767) );
  XOR2_X1 U858 ( .A(KEYINPUT34), .B(KEYINPUT89), .Z(n766) );
  XNOR2_X1 U859 ( .A(n767), .B(n766), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n894), .A2(G116), .ZN(n768) );
  XNOR2_X1 U861 ( .A(n768), .B(KEYINPUT90), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G128), .A2(n895), .ZN(n769) );
  NAND2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n771), .Z(n772) );
  NOR2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U866 ( .A(n774), .B(KEYINPUT36), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n776), .B(n775), .ZN(n883) );
  XNOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .ZN(n827) );
  NOR2_X1 U869 ( .A1(n883), .A2(n827), .ZN(n995) );
  NAND2_X1 U870 ( .A1(n829), .A2(n995), .ZN(n825) );
  NAND2_X1 U871 ( .A1(n894), .A2(G117), .ZN(n777) );
  XOR2_X1 U872 ( .A(KEYINPUT93), .B(n777), .Z(n779) );
  NAND2_X1 U873 ( .A1(n895), .A2(G129), .ZN(n778) );
  NAND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U875 ( .A(KEYINPUT94), .B(n780), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n898), .A2(G105), .ZN(n781) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n900), .A2(G141), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n885) );
  NAND2_X1 U881 ( .A1(n885), .A2(G1996), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G95), .A2(n898), .ZN(n787) );
  NAND2_X1 U883 ( .A1(G107), .A2(n894), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U885 ( .A1(G131), .A2(n900), .ZN(n789) );
  NAND2_X1 U886 ( .A1(G119), .A2(n895), .ZN(n788) );
  NAND2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n891) );
  NAND2_X1 U889 ( .A1(G1991), .A2(n891), .ZN(n792) );
  NAND2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U891 ( .A(n794), .B(KEYINPUT95), .ZN(n1003) );
  INV_X1 U892 ( .A(n1003), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n795), .A2(n829), .ZN(n819) );
  NAND2_X1 U894 ( .A1(n825), .A2(n819), .ZN(n812) );
  INV_X1 U895 ( .A(n812), .ZN(n796) );
  AND2_X1 U896 ( .A1(n933), .A2(n796), .ZN(n797) );
  NAND2_X1 U897 ( .A1(n798), .A2(n797), .ZN(n814) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n803) );
  NOR2_X1 U899 ( .A1(G2090), .A2(G303), .ZN(n801) );
  NAND2_X1 U900 ( .A1(G8), .A2(n801), .ZN(n802) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U902 ( .A1(n804), .A2(n807), .ZN(n810) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n805) );
  XOR2_X1 U904 ( .A(n805), .B(KEYINPUT24), .Z(n806) );
  NOR2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U906 ( .A(KEYINPUT97), .B(n808), .Z(n809) );
  NOR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n816), .B(n815), .ZN(n818) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n931) );
  NAND2_X1 U912 ( .A1(n931), .A2(n829), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n832) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n885), .ZN(n998) );
  INV_X1 U915 ( .A(n819), .ZN(n822) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n891), .ZN(n991) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n991), .A2(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n998), .A2(n823), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n824), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n883), .A2(n827), .ZN(n1005) );
  NAND2_X1 U924 ( .A1(n828), .A2(n1005), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n917), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U930 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U933 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U938 ( .A(G286), .B(G301), .Z(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n843), .B(n938), .Z(n844) );
  NOR2_X1 U941 ( .A1(G37), .A2(n844), .ZN(G397) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2678), .B(KEYINPUT108), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT107), .B(G2072), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2090), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(G2096), .B(G2100), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U951 ( .A(G2078), .B(G2084), .Z(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1966), .B(G1971), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1976), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(n857), .B(KEYINPUT41), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n864) );
  XOR2_X1 U959 ( .A(G2474), .B(G1956), .Z(n862) );
  XOR2_X1 U960 ( .A(G1981), .B(n860), .Z(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G112), .A2(n894), .ZN(n871) );
  NAND2_X1 U964 ( .A1(G100), .A2(n898), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G136), .A2(n900), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n895), .A2(G124), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT44), .B(n867), .Z(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT109), .ZN(G162) );
  XOR2_X1 U972 ( .A(n990), .B(G162), .Z(n874) );
  XNOR2_X1 U973 ( .A(G164), .B(G160), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n887) );
  NAND2_X1 U975 ( .A1(G103), .A2(n898), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G139), .A2(n900), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT113), .B(n877), .Z(n882) );
  NAND2_X1 U979 ( .A1(G115), .A2(n894), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G127), .A2(n895), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n1007) );
  XOR2_X1 U984 ( .A(n883), .B(n1007), .Z(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n893) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(KEYINPUT114), .Z(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n908) );
  NAND2_X1 U992 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n906) );
  NAND2_X1 U995 ( .A1(n898), .A2(G106), .ZN(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT110), .B(n899), .ZN(n903) );
  NAND2_X1 U997 ( .A1(n900), .A2(G142), .ZN(n901) );
  XOR2_X1 U998 ( .A(KEYINPUT111), .B(n901), .Z(n902) );
  NAND2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n904), .B(KEYINPUT45), .Z(n905) );
  NOR2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n911), .ZN(n915) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n916), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(KEYINPUT115), .B(n912), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(n913), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n916), .ZN(G319) );
  INV_X1 U1013 ( .A(n917), .ZN(G223) );
  XNOR2_X1 U1014 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1022) );
  XOR2_X1 U1015 ( .A(G1956), .B(KEYINPUT121), .Z(n918) );
  XOR2_X1 U1016 ( .A(n918), .B(G299), .Z(n920) );
  NAND2_X1 U1017 ( .A1(G1971), .A2(G303), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n929) );
  XOR2_X1 U1021 ( .A(G171), .B(G1961), .Z(n927) );
  XOR2_X1 U1022 ( .A(n925), .B(G1348), .Z(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(KEYINPUT122), .B(n932), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(G168), .B(G1966), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(n935), .B(KEYINPUT57), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(G1341), .B(n938), .ZN(n939) );
  NOR2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n942) );
  XOR2_X1 U1033 ( .A(G16), .B(KEYINPUT56), .Z(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n1020) );
  XOR2_X1 U1035 ( .A(G5), .B(G1961), .Z(n956) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G21), .ZN(n954) );
  XNOR2_X1 U1037 ( .A(G1981), .B(G6), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(KEYINPUT59), .B(G4), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(KEYINPUT123), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(G1348), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G1956), .B(G20), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT60), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT124), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(G1976), .B(G23), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G1971), .B(G22), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G1986), .B(G24), .Z(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT125), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(G11), .ZN(n989) );
  XOR2_X1 U1061 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1014) );
  XOR2_X1 U1062 ( .A(G1991), .B(G25), .Z(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(G28), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(G1996), .B(G32), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G2067), .B(G26), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G27), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1072 ( .A(KEYINPUT53), .B(n978), .Z(n981) );
  XOR2_X1 U1073 ( .A(G34), .B(KEYINPUT54), .Z(n979) );
  XNOR2_X1 U1074 ( .A(G2084), .B(n979), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1076 ( .A(KEYINPUT119), .B(G2090), .Z(n982) );
  XNOR2_X1 U1077 ( .A(G35), .B(n982), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n1014), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n986), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT120), .B(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n1018) );
  XNOR2_X1 U1083 ( .A(G160), .B(G2084), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT116), .B(n996), .Z(n1001) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT51), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT117), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1007), .Z(n1009) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1010), .Z(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1022), .B(n1021), .ZN(G311) );
  XNOR2_X1 U1106 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

