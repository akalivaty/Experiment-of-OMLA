

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742;

  BUF_X1 U378 ( .A(n567), .Z(n589) );
  INV_X2 U379 ( .A(G953), .ZN(n731) );
  NOR2_X1 U380 ( .A1(n738), .A2(n742), .ZN(n521) );
  AND2_X2 U381 ( .A1(n543), .A2(n381), .ZN(n380) );
  NOR2_X1 U382 ( .A1(n619), .A2(n600), .ZN(n465) );
  XNOR2_X2 U383 ( .A(n465), .B(n464), .ZN(n524) );
  NOR2_X1 U384 ( .A1(n741), .A2(n636), .ZN(n582) );
  NOR2_X1 U385 ( .A1(n658), .A2(n656), .ZN(n519) );
  AND2_X2 U386 ( .A1(n690), .A2(n422), .ZN(n705) );
  NOR2_X1 U387 ( .A1(n594), .A2(n572), .ZN(n574) );
  XNOR2_X1 U388 ( .A(n519), .B(n518), .ZN(n695) );
  NOR2_X1 U389 ( .A1(n560), .A2(n569), .ZN(n366) );
  XNOR2_X1 U390 ( .A(n410), .B(KEYINPUT102), .ZN(n560) );
  OR2_X2 U391 ( .A1(n668), .A2(n667), .ZN(n410) );
  XNOR2_X1 U392 ( .A(n603), .B(KEYINPUT111), .ZN(n604) );
  XNOR2_X1 U393 ( .A(n401), .B(n400), .ZN(n715) );
  XOR2_X1 U394 ( .A(n485), .B(n495), .Z(n727) );
  NAND2_X1 U395 ( .A1(n600), .A2(KEYINPUT2), .ZN(n419) );
  XNOR2_X1 U396 ( .A(n428), .B(n427), .ZN(n467) );
  XNOR2_X1 U397 ( .A(n460), .B(n461), .ZN(n428) );
  XNOR2_X1 U398 ( .A(n457), .B(G110), .ZN(n484) );
  XNOR2_X1 U399 ( .A(n730), .B(KEYINPUT74), .ZN(n361) );
  BUF_X1 U400 ( .A(n694), .Z(n354) );
  BUF_X1 U401 ( .A(n690), .Z(n355) );
  XNOR2_X1 U402 ( .A(n366), .B(n562), .ZN(n694) );
  XNOR2_X1 U403 ( .A(n408), .B(n363), .ZN(n712) );
  NOR2_X1 U404 ( .A1(n694), .A2(n589), .ZN(n563) );
  NAND2_X1 U405 ( .A1(n597), .A2(KEYINPUT86), .ZN(n389) );
  NAND2_X1 U406 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U407 ( .A1(n585), .A2(KEYINPUT44), .ZN(n593) );
  XOR2_X1 U408 ( .A(G131), .B(G140), .Z(n485) );
  OR2_X1 U409 ( .A1(G237), .A2(G902), .ZN(n466) );
  XNOR2_X1 U410 ( .A(n455), .B(n387), .ZN(n495) );
  INV_X1 U411 ( .A(KEYINPUT10), .ZN(n387) );
  NOR2_X1 U412 ( .A1(G953), .A2(G237), .ZN(n469) );
  XNOR2_X1 U413 ( .A(n484), .B(n458), .ZN(n400) );
  XNOR2_X1 U414 ( .A(n467), .B(n459), .ZN(n401) );
  XOR2_X1 U415 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n458) );
  XOR2_X1 U416 ( .A(KEYINPUT82), .B(n544), .Z(n545) );
  NAND2_X1 U417 ( .A1(n582), .A2(n739), .ZN(n579) );
  NOR2_X1 U418 ( .A1(n391), .A2(n388), .ZN(n369) );
  NAND2_X1 U419 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U420 ( .A(n468), .B(n426), .ZN(n425) );
  INV_X1 U421 ( .A(G116), .ZN(n426) );
  XOR2_X1 U422 ( .A(KEYINPUT5), .B(G131), .Z(n468) );
  XNOR2_X1 U423 ( .A(G137), .B(G134), .ZN(n471) );
  XNOR2_X1 U424 ( .A(G101), .B(KEYINPUT70), .ZN(n427) );
  XNOR2_X1 U425 ( .A(n433), .B(n409), .ZN(n500) );
  XNOR2_X1 U426 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n433) );
  NAND2_X1 U427 ( .A1(n731), .A2(G234), .ZN(n409) );
  INV_X1 U428 ( .A(n485), .ZN(n413) );
  XNOR2_X1 U429 ( .A(n487), .B(n486), .ZN(n488) );
  INV_X1 U430 ( .A(KEYINPUT77), .ZN(n486) );
  XNOR2_X1 U431 ( .A(G101), .B(G107), .ZN(n487) );
  XNOR2_X1 U432 ( .A(G104), .B(KEYINPUT91), .ZN(n457) );
  INV_X1 U433 ( .A(KEYINPUT48), .ZN(n405) );
  NOR2_X1 U434 ( .A1(n569), .A2(n424), .ZN(n423) );
  XNOR2_X1 U435 ( .A(n530), .B(n529), .ZN(n668) );
  XNOR2_X1 U436 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U437 ( .A(n474), .B(n417), .ZN(n671) );
  INV_X1 U438 ( .A(G472), .ZN(n417) );
  XNOR2_X1 U439 ( .A(n559), .B(KEYINPUT0), .ZN(n567) );
  BUF_X1 U440 ( .A(n671), .Z(n376) );
  NOR2_X1 U441 ( .A1(n712), .A2(G902), .ZN(n407) );
  XNOR2_X1 U442 ( .A(G140), .B(KEYINPUT94), .ZN(n501) );
  XNOR2_X1 U443 ( .A(G119), .B(G137), .ZN(n496) );
  XOR2_X1 U444 ( .A(G110), .B(G128), .Z(n497) );
  XNOR2_X1 U445 ( .A(G116), .B(G107), .ZN(n430) );
  XNOR2_X1 U446 ( .A(n445), .B(n360), .ZN(n446) );
  XNOR2_X1 U447 ( .A(KEYINPUT6), .B(n671), .ZN(n569) );
  BUF_X1 U448 ( .A(n668), .Z(n378) );
  XNOR2_X1 U449 ( .A(n368), .B(KEYINPUT22), .ZN(n575) );
  NOR2_X1 U450 ( .A1(n567), .A2(n402), .ZN(n368) );
  NAND2_X1 U451 ( .A1(n403), .A2(n568), .ZN(n402) );
  INV_X1 U452 ( .A(n656), .ZN(n403) );
  NOR2_X1 U453 ( .A1(n545), .A2(n357), .ZN(n381) );
  INV_X1 U454 ( .A(KEYINPUT72), .ZN(n578) );
  XNOR2_X1 U455 ( .A(n550), .B(n372), .ZN(n517) );
  INV_X1 U456 ( .A(KEYINPUT38), .ZN(n372) );
  XNOR2_X1 U457 ( .A(n467), .B(n377), .ZN(n473) );
  XNOR2_X1 U458 ( .A(n425), .B(n470), .ZN(n377) );
  XNOR2_X1 U459 ( .A(n490), .B(n411), .ZN(n699) );
  XNOR2_X1 U460 ( .A(n414), .B(n412), .ZN(n411) );
  XNOR2_X1 U461 ( .A(n488), .B(n413), .ZN(n412) );
  XNOR2_X1 U462 ( .A(n456), .B(n399), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n453), .B(KEYINPUT18), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n421), .B(KEYINPUT75), .ZN(n690) );
  NAND2_X1 U465 ( .A1(n386), .A2(n423), .ZN(n546) );
  INV_X1 U466 ( .A(n374), .ZN(n386) );
  INV_X1 U467 ( .A(n410), .ZN(n586) );
  NAND2_X1 U468 ( .A1(n524), .A2(n652), .ZN(n365) );
  XNOR2_X1 U469 ( .A(n531), .B(n532), .ZN(n643) );
  XNOR2_X1 U470 ( .A(n504), .B(n499), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n435), .B(n375), .ZN(n707) );
  XNOR2_X1 U472 ( .A(n434), .B(n436), .ZN(n375) );
  XNOR2_X1 U473 ( .A(n611), .B(n610), .ZN(n612) );
  AND2_X1 U474 ( .A1(n575), .A2(n416), .ZN(n576) );
  BUF_X1 U475 ( .A(n643), .Z(n374) );
  NAND2_X1 U476 ( .A1(n590), .A2(n416), .ZN(n631) );
  OR2_X1 U477 ( .A1(n594), .A2(n663), .ZN(n595) );
  AND2_X1 U478 ( .A1(n423), .A2(n524), .ZN(n356) );
  AND2_X1 U479 ( .A1(n528), .A2(n527), .ZN(n357) );
  XOR2_X1 U480 ( .A(KEYINPUT25), .B(n494), .Z(n358) );
  XOR2_X1 U481 ( .A(KEYINPUT69), .B(G469), .Z(n359) );
  AND2_X1 U482 ( .A1(G214), .A2(n469), .ZN(n360) );
  AND2_X1 U483 ( .A1(n533), .A2(n652), .ZN(n362) );
  XOR2_X1 U484 ( .A(n498), .B(n503), .Z(n363) );
  INV_X1 U485 ( .A(n524), .ZN(n550) );
  INV_X2 U486 ( .A(G146), .ZN(n415) );
  XNOR2_X1 U487 ( .A(KEYINPUT15), .B(G902), .ZN(n491) );
  XNOR2_X1 U488 ( .A(n715), .B(n397), .ZN(n619) );
  XOR2_X1 U489 ( .A(n598), .B(KEYINPUT45), .Z(n364) );
  NAND2_X1 U490 ( .A1(n575), .A2(n569), .ZN(n594) );
  NOR2_X2 U491 ( .A1(n596), .A2(n595), .ZN(n628) );
  XNOR2_X2 U492 ( .A(n365), .B(KEYINPUT19), .ZN(n558) );
  XNOR2_X2 U493 ( .A(n566), .B(KEYINPUT35), .ZN(n585) );
  NAND2_X1 U494 ( .A1(n705), .A2(G472), .ZN(n605) );
  NAND2_X1 U495 ( .A1(n705), .A2(G210), .ZN(n623) );
  NAND2_X1 U496 ( .A1(n705), .A2(G475), .ZN(n613) );
  XNOR2_X1 U497 ( .A(n367), .B(n405), .ZN(n404) );
  NAND2_X1 U498 ( .A1(n406), .A2(n379), .ZN(n367) );
  XNOR2_X1 U499 ( .A(n512), .B(n429), .ZN(n738) );
  XOR2_X1 U500 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n502) );
  NOR2_X2 U501 ( .A1(n588), .A2(n513), .ZN(n508) );
  NOR2_X2 U502 ( .A1(n538), .A2(n517), .ZN(n371) );
  XNOR2_X1 U503 ( .A(n371), .B(KEYINPUT39), .ZN(n552) );
  NAND2_X1 U504 ( .A1(n581), .A2(n580), .ZN(n396) );
  NAND2_X1 U505 ( .A1(n369), .A2(n396), .ZN(n395) );
  XNOR2_X2 U506 ( .A(n370), .B(n359), .ZN(n530) );
  OR2_X2 U507 ( .A1(n699), .A2(G902), .ZN(n370) );
  XNOR2_X2 U508 ( .A(n472), .B(n471), .ZN(n729) );
  XNOR2_X2 U509 ( .A(n451), .B(n452), .ZN(n472) );
  XNOR2_X2 U510 ( .A(KEYINPUT20), .B(n492), .ZN(n505) );
  XNOR2_X1 U511 ( .A(n520), .B(KEYINPUT42), .ZN(n742) );
  NAND2_X1 U512 ( .A1(n383), .A2(n373), .ZN(n534) );
  NAND2_X1 U513 ( .A1(n385), .A2(n356), .ZN(n373) );
  NOR2_X2 U514 ( .A1(n687), .A2(n599), .ZN(n421) );
  XNOR2_X1 U515 ( .A(n489), .B(n484), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n380), .B(KEYINPUT68), .ZN(n379) );
  NAND2_X1 U517 ( .A1(n382), .A2(n356), .ZN(n384) );
  INV_X1 U518 ( .A(n643), .ZN(n382) );
  NAND2_X1 U519 ( .A1(n384), .A2(KEYINPUT36), .ZN(n383) );
  NOR2_X1 U520 ( .A1(n643), .A2(KEYINPUT36), .ZN(n385) );
  XNOR2_X2 U521 ( .A(n415), .B(G125), .ZN(n455) );
  NAND2_X1 U522 ( .A1(n628), .A2(KEYINPUT86), .ZN(n390) );
  NAND2_X1 U523 ( .A1(n392), .A2(n584), .ZN(n391) );
  NAND2_X1 U524 ( .A1(n394), .A2(n393), .ZN(n392) );
  INV_X1 U525 ( .A(n628), .ZN(n393) );
  NOR2_X1 U526 ( .A1(n597), .A2(KEYINPUT86), .ZN(n394) );
  XNOR2_X2 U527 ( .A(n395), .B(n364), .ZN(n687) );
  INV_X1 U528 ( .A(n452), .ZN(n450) );
  XNOR2_X2 U529 ( .A(G128), .B(G143), .ZN(n452) );
  XNOR2_X1 U530 ( .A(n472), .B(n398), .ZN(n397) );
  NAND2_X1 U531 ( .A1(n404), .A2(n651), .ZN(n601) );
  XNOR2_X1 U532 ( .A(n521), .B(KEYINPUT46), .ZN(n406) );
  XNOR2_X2 U533 ( .A(n407), .B(n358), .ZN(n570) );
  NOR2_X2 U534 ( .A1(n378), .A2(n534), .ZN(n648) );
  XNOR2_X2 U535 ( .A(n729), .B(n415), .ZN(n490) );
  INV_X1 U536 ( .A(n376), .ZN(n416) );
  NAND2_X1 U537 ( .A1(n418), .A2(n361), .ZN(n420) );
  NOR2_X1 U538 ( .A1(n687), .A2(n491), .ZN(n418) );
  NAND2_X1 U539 ( .A1(n420), .A2(n419), .ZN(n422) );
  NAND2_X1 U540 ( .A1(n522), .A2(n536), .ZN(n531) );
  NAND2_X1 U541 ( .A1(n663), .A2(n362), .ZN(n424) );
  OR2_X2 U542 ( .A1(n601), .A2(n554), .ZN(n599) );
  XNOR2_X1 U543 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X2 U544 ( .A(G113), .B(KEYINPUT3), .ZN(n460) );
  XNOR2_X1 U545 ( .A(n490), .B(n473), .ZN(n602) );
  XNOR2_X2 U546 ( .A(n449), .B(n448), .ZN(n537) );
  NOR2_X2 U547 ( .A1(G902), .A2(n609), .ZN(n449) );
  XOR2_X1 U548 ( .A(n511), .B(KEYINPUT108), .Z(n429) );
  INV_X1 U549 ( .A(KEYINPUT85), .ZN(n535) );
  XNOR2_X1 U550 ( .A(n579), .B(n578), .ZN(n581) );
  INV_X1 U551 ( .A(KEYINPUT11), .ZN(n441) );
  XNOR2_X1 U552 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U554 ( .A(KEYINPUT30), .ZN(n476) );
  INV_X1 U555 ( .A(KEYINPUT93), .ZN(n462) );
  XNOR2_X1 U556 ( .A(n447), .B(G475), .ZN(n448) );
  XNOR2_X1 U557 ( .A(n561), .B(KEYINPUT71), .ZN(n562) );
  XNOR2_X1 U558 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n529) );
  NOR2_X2 U559 ( .A1(n601), .A2(n650), .ZN(n730) );
  XNOR2_X1 U560 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U561 ( .A(n709), .B(n708), .ZN(n710) );
  INV_X1 U562 ( .A(n491), .ZN(n600) );
  XNOR2_X1 U563 ( .A(n430), .B(G122), .ZN(n459) );
  XNOR2_X1 U564 ( .A(n450), .B(KEYINPUT9), .ZN(n431) );
  XNOR2_X1 U565 ( .A(n431), .B(KEYINPUT99), .ZN(n432) );
  XOR2_X1 U566 ( .A(n459), .B(n432), .Z(n435) );
  NAND2_X1 U567 ( .A1(G217), .A2(n500), .ZN(n434) );
  XOR2_X1 U568 ( .A(G134), .B(KEYINPUT7), .Z(n436) );
  NOR2_X1 U569 ( .A1(G902), .A2(n707), .ZN(n438) );
  XNOR2_X1 U570 ( .A(KEYINPUT100), .B(G478), .ZN(n437) );
  XNOR2_X1 U571 ( .A(n438), .B(n437), .ZN(n536) );
  XOR2_X1 U572 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n440) );
  XNOR2_X1 U573 ( .A(G143), .B(G104), .ZN(n439) );
  XNOR2_X1 U574 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U575 ( .A(G113), .B(G122), .ZN(n442) );
  XNOR2_X1 U576 ( .A(n446), .B(n727), .ZN(n609) );
  XNOR2_X1 U577 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n447) );
  XOR2_X1 U578 ( .A(n537), .B(KEYINPUT98), .Z(n522) );
  XNOR2_X1 U579 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n451) );
  NAND2_X1 U580 ( .A1(n731), .A2(G224), .ZN(n453) );
  XOR2_X1 U581 ( .A(KEYINPUT78), .B(KEYINPUT17), .Z(n454) );
  XNOR2_X2 U582 ( .A(G119), .B(KEYINPUT92), .ZN(n461) );
  NAND2_X1 U583 ( .A1(G210), .A2(n466), .ZN(n463) );
  NAND2_X1 U584 ( .A1(G214), .A2(n466), .ZN(n652) );
  NAND2_X1 U585 ( .A1(n469), .A2(G210), .ZN(n470) );
  NOR2_X1 U586 ( .A1(n602), .A2(G902), .ZN(n474) );
  NAND2_X1 U587 ( .A1(n652), .A2(n671), .ZN(n475) );
  XNOR2_X1 U588 ( .A(n475), .B(KEYINPUT106), .ZN(n477) );
  XNOR2_X1 U589 ( .A(n477), .B(n476), .ZN(n510) );
  NAND2_X1 U590 ( .A1(G234), .A2(G237), .ZN(n478) );
  XNOR2_X1 U591 ( .A(n478), .B(KEYINPUT14), .ZN(n683) );
  OR2_X1 U592 ( .A1(n731), .A2(G902), .ZN(n479) );
  NAND2_X1 U593 ( .A1(n683), .A2(n479), .ZN(n481) );
  NOR2_X1 U594 ( .A1(G953), .A2(G952), .ZN(n480) );
  NOR2_X1 U595 ( .A1(n481), .A2(n480), .ZN(n556) );
  NAND2_X1 U596 ( .A1(G953), .A2(G900), .ZN(n482) );
  NAND2_X1 U597 ( .A1(n556), .A2(n482), .ZN(n483) );
  XOR2_X1 U598 ( .A(KEYINPUT79), .B(n483), .Z(n513) );
  NAND2_X1 U599 ( .A1(G227), .A2(n731), .ZN(n489) );
  NAND2_X1 U600 ( .A1(G234), .A2(n491), .ZN(n492) );
  NAND2_X1 U601 ( .A1(n505), .A2(G217), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n493), .B(KEYINPUT95), .ZN(n494) );
  INV_X1 U603 ( .A(n495), .ZN(n499) );
  XNOR2_X1 U604 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U605 ( .A1(n500), .A2(G221), .ZN(n504) );
  XNOR2_X1 U606 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U607 ( .A1(n505), .A2(G221), .ZN(n506) );
  XOR2_X1 U608 ( .A(n506), .B(KEYINPUT21), .Z(n568) );
  NAND2_X1 U609 ( .A1(n570), .A2(n568), .ZN(n667) );
  INV_X1 U610 ( .A(n667), .ZN(n507) );
  NAND2_X1 U611 ( .A1(n530), .A2(n507), .ZN(n588) );
  XNOR2_X1 U612 ( .A(KEYINPUT76), .B(n508), .ZN(n509) );
  NAND2_X1 U613 ( .A1(n510), .A2(n509), .ZN(n538) );
  NOR2_X1 U614 ( .A1(n531), .A2(n552), .ZN(n512) );
  XNOR2_X1 U615 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n511) );
  INV_X1 U616 ( .A(n568), .ZN(n664) );
  NOR2_X1 U617 ( .A1(n664), .A2(n513), .ZN(n533) );
  NAND2_X1 U618 ( .A1(n671), .A2(n533), .ZN(n514) );
  NOR2_X1 U619 ( .A1(n570), .A2(n514), .ZN(n515) );
  XNOR2_X1 U620 ( .A(KEYINPUT28), .B(n515), .ZN(n516) );
  NAND2_X1 U621 ( .A1(n516), .A2(n530), .ZN(n523) );
  INV_X1 U622 ( .A(n517), .ZN(n653) );
  NAND2_X1 U623 ( .A1(n653), .A2(n652), .ZN(n658) );
  NAND2_X1 U624 ( .A1(n536), .A2(n537), .ZN(n656) );
  XNOR2_X1 U625 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n518) );
  NOR2_X1 U626 ( .A1(n523), .A2(n695), .ZN(n520) );
  OR2_X1 U627 ( .A1(n522), .A2(n536), .ZN(n646) );
  NAND2_X1 U628 ( .A1(n531), .A2(n646), .ZN(n657) );
  XOR2_X1 U629 ( .A(KEYINPUT47), .B(n657), .Z(n528) );
  INV_X1 U630 ( .A(KEYINPUT47), .ZN(n526) );
  INV_X1 U631 ( .A(n523), .ZN(n525) );
  NAND2_X1 U632 ( .A1(n525), .A2(n558), .ZN(n640) );
  NAND2_X1 U633 ( .A1(n526), .A2(n640), .ZN(n527) );
  INV_X1 U634 ( .A(n570), .ZN(n663) );
  INV_X1 U635 ( .A(KEYINPUT103), .ZN(n532) );
  XNOR2_X1 U636 ( .A(n648), .B(n535), .ZN(n542) );
  NOR2_X1 U637 ( .A1(n537), .A2(n536), .ZN(n564) );
  INV_X1 U638 ( .A(n564), .ZN(n541) );
  NOR2_X1 U639 ( .A1(n550), .A2(n538), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n539), .B(KEYINPUT107), .ZN(n540) );
  NOR2_X1 U641 ( .A1(n541), .A2(n540), .ZN(n639) );
  NOR2_X1 U642 ( .A1(n542), .A2(n639), .ZN(n543) );
  NAND2_X1 U643 ( .A1(n640), .A2(KEYINPUT47), .ZN(n544) );
  INV_X1 U644 ( .A(n378), .ZN(n596) );
  XNOR2_X1 U645 ( .A(KEYINPUT104), .B(n546), .ZN(n547) );
  NOR2_X1 U646 ( .A1(n596), .A2(n547), .ZN(n548) );
  XNOR2_X1 U647 ( .A(KEYINPUT43), .B(n548), .ZN(n549) );
  XNOR2_X1 U648 ( .A(n549), .B(KEYINPUT105), .ZN(n551) );
  NAND2_X1 U649 ( .A1(n551), .A2(n550), .ZN(n651) );
  INV_X1 U650 ( .A(KEYINPUT2), .ZN(n688) );
  NOR2_X1 U651 ( .A1(n646), .A2(n552), .ZN(n650) );
  OR2_X1 U652 ( .A1(n688), .A2(n650), .ZN(n553) );
  XNOR2_X1 U653 ( .A(KEYINPUT80), .B(n553), .ZN(n554) );
  NAND2_X1 U654 ( .A1(G898), .A2(G953), .ZN(n555) );
  AND2_X1 U655 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U656 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U657 ( .A(KEYINPUT33), .ZN(n561) );
  XNOR2_X1 U658 ( .A(n563), .B(KEYINPUT34), .ZN(n565) );
  NAND2_X1 U659 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U660 ( .A(n585), .ZN(n739) );
  NOR2_X1 U661 ( .A1(n378), .A2(n570), .ZN(n571) );
  XNOR2_X1 U662 ( .A(KEYINPUT101), .B(n571), .ZN(n572) );
  XNOR2_X1 U663 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n573) );
  XNOR2_X1 U664 ( .A(n574), .B(n573), .ZN(n741) );
  NAND2_X1 U665 ( .A1(n663), .A2(n576), .ZN(n577) );
  NOR2_X1 U666 ( .A1(n596), .A2(n577), .ZN(n636) );
  INV_X1 U667 ( .A(KEYINPUT44), .ZN(n580) );
  NAND2_X1 U668 ( .A1(KEYINPUT72), .A2(n582), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n583), .A2(KEYINPUT44), .ZN(n584) );
  NAND2_X1 U670 ( .A1(n376), .A2(n586), .ZN(n676) );
  NOR2_X1 U671 ( .A1(n589), .A2(n676), .ZN(n587) );
  XNOR2_X1 U672 ( .A(KEYINPUT31), .B(n587), .ZN(n645) );
  NOR2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n645), .A2(n631), .ZN(n591) );
  NAND2_X1 U675 ( .A1(n591), .A2(n657), .ZN(n592) );
  XNOR2_X1 U676 ( .A(KEYINPUT84), .B(KEYINPUT64), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT62), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n605), .B(n604), .ZN(n607) );
  NOR2_X1 U679 ( .A1(G952), .A2(n731), .ZN(n606) );
  XNOR2_X1 U680 ( .A(KEYINPUT90), .B(n606), .ZN(n714) );
  INV_X1 U681 ( .A(n714), .ZN(n624) );
  NAND2_X1 U682 ( .A1(n607), .A2(n624), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U684 ( .A(KEYINPUT89), .B(KEYINPUT120), .Z(n611) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT59), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(n624), .ZN(n616) );
  INV_X1 U688 ( .A(KEYINPUT60), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(G60) );
  XNOR2_X1 U690 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT81), .ZN(n618) );
  XNOR2_X1 U692 ( .A(KEYINPUT54), .B(n618), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT55), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n627) );
  INV_X1 U697 ( .A(KEYINPUT56), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(G51) );
  XOR2_X1 U699 ( .A(G101), .B(n628), .Z(n629) );
  XNOR2_X1 U700 ( .A(KEYINPUT112), .B(n629), .ZN(G3) );
  NOR2_X1 U701 ( .A1(n374), .A2(n631), .ZN(n630) );
  XOR2_X1 U702 ( .A(G104), .B(n630), .Z(G6) );
  NOR2_X1 U703 ( .A1(n631), .A2(n646), .ZN(n635) );
  XOR2_X1 U704 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n633) );
  XNOR2_X1 U705 ( .A(G107), .B(KEYINPUT26), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(G9) );
  XOR2_X1 U708 ( .A(n636), .B(G110), .Z(G12) );
  NOR2_X1 U709 ( .A1(n640), .A2(n646), .ZN(n638) );
  XNOR2_X1 U710 ( .A(G128), .B(KEYINPUT29), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G30) );
  XOR2_X1 U712 ( .A(G143), .B(n639), .Z(G45) );
  NOR2_X1 U713 ( .A1(n374), .A2(n640), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT114), .B(n641), .Z(n642) );
  XNOR2_X1 U715 ( .A(G146), .B(n642), .ZN(G48) );
  NOR2_X1 U716 ( .A1(n374), .A2(n645), .ZN(n644) );
  XOR2_X1 U717 ( .A(G113), .B(n644), .Z(G15) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U719 ( .A(G116), .B(n647), .Z(G18) );
  XNOR2_X1 U720 ( .A(G125), .B(n648), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n649), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U722 ( .A(G134), .B(n650), .Z(G36) );
  XNOR2_X1 U723 ( .A(G140), .B(n651), .ZN(G42) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U725 ( .A(KEYINPUT117), .B(n654), .Z(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n661) );
  INV_X1 U727 ( .A(n657), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n354), .A2(n662), .ZN(n680) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n665), .B(KEYINPUT115), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT49), .B(n666), .ZN(n674) );
  XOR2_X1 U734 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n670) );
  NAND2_X1 U735 ( .A1(n378), .A2(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n670), .B(n669), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n672), .A2(n376), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(KEYINPUT51), .B(n677), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n695), .A2(n678), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  XNOR2_X1 U744 ( .A(n682), .B(KEYINPUT118), .ZN(n685) );
  NAND2_X1 U745 ( .A1(G952), .A2(n683), .ZN(n684) );
  NOR2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U747 ( .A1(G953), .A2(n686), .ZN(n693) );
  INV_X1 U748 ( .A(n687), .ZN(n718) );
  NAND2_X1 U749 ( .A1(n718), .A2(n730), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U751 ( .A1(n691), .A2(n355), .ZN(n692) );
  NAND2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U753 ( .A1(n695), .A2(n354), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U755 ( .A(KEYINPUT53), .B(n698), .ZN(G75) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n701) );
  XNOR2_X1 U757 ( .A(n699), .B(KEYINPUT119), .ZN(n700) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U759 ( .A1(n705), .A2(G469), .ZN(n702) );
  XOR2_X1 U760 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U761 ( .A1(n714), .A2(n704), .ZN(G54) );
  NAND2_X1 U762 ( .A1(n705), .A2(G478), .ZN(n709) );
  XOR2_X1 U763 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n706) );
  NOR2_X1 U764 ( .A1(n714), .A2(n710), .ZN(G63) );
  NAND2_X1 U765 ( .A1(G217), .A2(n705), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U768 ( .A(KEYINPUT125), .B(n715), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n731), .A2(G898), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n717), .A2(n716), .ZN(n726) );
  NAND2_X1 U771 ( .A1(n718), .A2(n731), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(KEYINPUT124), .ZN(n724) );
  XOR2_X1 U773 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n721) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U775 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U776 ( .A1(n722), .A2(G898), .ZN(n723) );
  NAND2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(G69) );
  XOR2_X1 U779 ( .A(n727), .B(KEYINPUT126), .Z(n728) );
  XOR2_X1 U780 ( .A(n729), .B(n728), .Z(n733) );
  XOR2_X1 U781 ( .A(n733), .B(n730), .Z(n732) );
  NAND2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n737) );
  XNOR2_X1 U783 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U785 ( .A1(G953), .A2(n735), .ZN(n736) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U787 ( .A(n738), .B(G131), .Z(G33) );
  XOR2_X1 U788 ( .A(G122), .B(n739), .Z(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U790 ( .A(G119), .B(n741), .Z(G21) );
  XOR2_X1 U791 ( .A(G137), .B(n742), .Z(G39) );
endmodule

