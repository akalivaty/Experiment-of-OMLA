//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n206), .A2(new_n207), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n211), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n224), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(G274), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n226), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n256), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n257), .B1(new_n261), .B2(new_n219), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G232), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT68), .A2(G107), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT68), .A2(G107), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(G1698), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n265), .B1(new_n269), .B2(new_n263), .C1(new_n270), .C2(new_n213), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n226), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n251), .B2(new_n252), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n262), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G200), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n226), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n227), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n227), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT15), .B(G87), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n227), .A2(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n289), .A2(new_n291), .B1(new_n227), .B2(new_n218), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n280), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n280), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G77), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT69), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n295), .A2(new_n227), .A3(G1), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n280), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(G77), .A4(new_n300), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n218), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n293), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT70), .B1(new_n278), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n293), .A2(new_n307), .A3(new_n308), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT70), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n311), .B(new_n312), .C1(new_n277), .C2(new_n276), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n276), .A2(G190), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n309), .B1(new_n276), .B2(G169), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n309), .B(KEYINPUT71), .C1(G169), .C2(new_n276), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n276), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT72), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n326), .B1(new_n218), .B2(new_n263), .C1(new_n270), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n275), .ZN(new_n329));
  INV_X1    g0129(.A(new_n257), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G226), .B2(new_n260), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G169), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(G179), .ZN(new_n335));
  INV_X1    g0135(.A(new_n289), .ZN(new_n336));
  INV_X1    g0136(.A(new_n291), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n285), .A2(new_n336), .B1(G150), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n208), .A2(G20), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n294), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n304), .A2(G50), .A3(new_n300), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G50), .B2(new_n297), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n334), .A2(new_n335), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(G200), .A2(new_n332), .B1(new_n343), .B2(KEYINPUT9), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n333), .A2(G190), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n343), .A2(KEYINPUT9), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT10), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT10), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n315), .A2(new_n322), .A3(KEYINPUT72), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n325), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n327), .A2(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G33), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n263), .A2(G226), .A3(G1698), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n263), .A2(KEYINPUT76), .A3(new_n356), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n275), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n275), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n299), .B1(G41), .B2(G45), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n253), .A2(G232), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n257), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n257), .B2(new_n372), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n374), .A2(new_n375), .A3(G190), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n366), .A2(new_n275), .ZN(new_n378));
  INV_X1    g0178(.A(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n257), .A2(new_n372), .A3(new_n373), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n277), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n336), .A2(new_n300), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(new_n298), .B1(new_n297), .B2(new_n336), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n357), .A2(new_n359), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(new_n227), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n202), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n263), .B2(G20), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n358), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT7), .B(new_n227), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(KEYINPUT75), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n291), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n398), .B(new_n400), .C1(new_n401), .C2(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n294), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n202), .B1(new_n392), .B2(new_n395), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n201), .A2(new_n202), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n206), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n400), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n398), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n386), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n383), .A2(new_n384), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n383), .A2(new_n410), .A3(new_n384), .A4(KEYINPUT17), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n392), .A2(KEYINPUT75), .A3(new_n395), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n392), .B2(KEYINPUT75), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n402), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n409), .A3(new_n280), .ZN(new_n418));
  INV_X1    g0218(.A(new_n386), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n374), .A2(new_n375), .ZN(new_n421));
  AOI21_X1  g0221(.A(G169), .B1(new_n421), .B2(new_n367), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n369), .A2(new_n320), .A3(new_n370), .A4(new_n421), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT18), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n420), .A2(new_n427), .A3(new_n423), .A4(new_n424), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n413), .A2(new_n414), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT80), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n263), .A2(G226), .A3(new_n264), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n275), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n330), .B1(G238), .B2(new_n260), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT13), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(G169), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT14), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n440), .A2(new_n444), .A3(G169), .A4(new_n441), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(KEYINPUT73), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT73), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n436), .A2(new_n437), .B1(new_n447), .B2(KEYINPUT13), .ZN(new_n448));
  OAI21_X1  g0248(.A(G179), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n443), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n303), .A2(new_n202), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT12), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n304), .A2(G68), .A3(new_n300), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n286), .A2(new_n218), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n291), .A2(new_n207), .B1(new_n227), .B2(G68), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n280), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT11), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n440), .A2(G200), .A3(new_n441), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G190), .B1(new_n446), .B2(new_n448), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n450), .A2(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n355), .A2(new_n430), .A3(new_n431), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n430), .A2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT80), .B1(new_n467), .B2(new_n354), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n294), .B(new_n297), .C1(G1), .C2(new_n290), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n220), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n296), .A2(G20), .A3(new_n220), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT25), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n220), .A2(G20), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  OAI22_X1  g0277(.A1(KEYINPUT23), .A2(new_n476), .B1(new_n281), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n266), .A2(G20), .A3(new_n267), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(KEYINPUT23), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n357), .A2(new_n359), .A3(new_n227), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n263), .A2(new_n483), .A3(new_n227), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n475), .B1(new_n491), .B2(new_n280), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n357), .A2(new_n359), .A3(G257), .A4(G1698), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n263), .A2(KEYINPUT88), .A3(G257), .A4(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n263), .A2(G250), .A3(new_n264), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n275), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n299), .A2(G45), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n221), .A3(new_n259), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n504), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n255), .A2(G1), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n253), .A3(G274), .A4(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n506), .B1(new_n500), .B2(new_n275), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n277), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n501), .A2(new_n512), .A3(new_n507), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n519));
  INV_X1    g0319(.A(G190), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT89), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(new_n521), .A3(new_n512), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n493), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n513), .A2(new_n521), .A3(new_n512), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n513), .B2(new_n512), .ZN(new_n526));
  OAI21_X1  g0326(.A(G169), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n509), .A2(G179), .A3(new_n512), .A4(new_n515), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n492), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n279), .A2(new_n226), .B1(G20), .B2(new_n477), .ZN(new_n531));
  AOI21_X1  g0331(.A(G20), .B1(G33), .B2(G283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n290), .A2(G97), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT84), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(KEYINPUT20), .B(new_n531), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n470), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G116), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n303), .A2(new_n477), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n510), .A2(new_n511), .B1(new_n251), .B2(new_n252), .ZN(new_n546));
  INV_X1    g0346(.A(G274), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n259), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(G270), .B1(new_n548), .B2(new_n505), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n357), .A2(new_n359), .A3(G257), .A4(new_n264), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n357), .A2(new_n359), .A3(G264), .A4(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(G303), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n263), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n275), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n545), .A2(KEYINPUT21), .A3(G169), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(G169), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n544), .B1(new_n470), .B2(new_n477), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n539), .B2(new_n540), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n549), .A2(new_n554), .A3(G179), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n545), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT85), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n277), .B1(new_n549), .B2(new_n554), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n545), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n555), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n560), .B(KEYINPUT85), .C1(new_n568), .C2(new_n277), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(G190), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT86), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(new_n569), .A3(new_n573), .A4(new_n570), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n564), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n357), .A2(new_n359), .A3(G244), .A4(new_n264), .ZN(new_n576));
  NOR2_X1   g0376(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n577), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n263), .A2(G244), .A3(new_n264), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G283), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n578), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n275), .ZN(new_n584));
  INV_X1    g0384(.A(new_n504), .ZN(new_n585));
  NOR2_X1   g0385(.A1(KEYINPUT5), .A2(G41), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n511), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G257), .A3(new_n253), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n512), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G179), .ZN(new_n592));
  INV_X1    g0392(.A(G97), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n303), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n470), .B2(new_n593), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n593), .A2(new_n220), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n220), .A2(KEYINPUT6), .A3(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(G20), .B1(G77), .B2(new_n337), .ZN(new_n602));
  INV_X1    g0402(.A(new_n395), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n268), .B1(new_n603), .B2(new_n388), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n595), .B1(new_n605), .B2(new_n280), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n589), .B1(new_n583), .B2(new_n275), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n592), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT82), .ZN(new_n611));
  AOI211_X1 g0411(.A(G190), .B(new_n589), .C1(new_n583), .C2(new_n275), .ZN(new_n612));
  AOI21_X1  g0412(.A(G200), .B1(new_n584), .B2(new_n590), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n606), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n584), .A2(new_n520), .A3(new_n590), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(G200), .B2(new_n607), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n611), .B1(new_n617), .B2(new_n606), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n610), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n227), .B1(new_n434), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n214), .A2(new_n593), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n268), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n263), .A2(new_n227), .A3(G68), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n593), .B1(new_n282), .B2(new_n284), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(KEYINPUT19), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n280), .B1(new_n303), .B2(new_n287), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n542), .A2(G87), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n357), .A2(new_n359), .A3(G244), .A4(G1698), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n357), .A2(new_n359), .A3(G238), .A4(new_n264), .ZN(new_n631));
  NAND2_X1  g0431(.A1(G33), .A2(G116), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n275), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n511), .A2(new_n215), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n548), .A2(new_n511), .B1(new_n253), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT83), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(new_n636), .A3(KEYINPUT83), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G190), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n640), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT83), .B1(new_n634), .B2(new_n636), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n629), .B(new_n641), .C1(new_n644), .C2(new_n277), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n639), .A2(new_n320), .A3(new_n640), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n627), .B1(new_n287), .B2(new_n470), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n646), .B(new_n647), .C1(new_n644), .C2(G169), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n619), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n469), .A2(new_n530), .A3(new_n575), .A4(new_n650), .ZN(G372));
  AOI21_X1  g0451(.A(new_n514), .B1(new_n501), .B2(new_n507), .ZN(new_n652));
  AOI211_X1 g0452(.A(KEYINPUT90), .B(new_n506), .C1(new_n500), .C2(new_n275), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(G200), .B1(new_n654), .B2(new_n512), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n525), .A2(new_n526), .A3(G190), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n492), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n606), .B1(new_n612), .B2(new_n613), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT82), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n609), .B1(new_n659), .B2(new_n614), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n637), .A2(G200), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n629), .A2(new_n641), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G169), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n637), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n646), .A2(new_n647), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n662), .A2(new_n665), .A3(KEYINPUT91), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT91), .B1(new_n662), .B2(new_n665), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n657), .B(new_n660), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n564), .ZN(new_n669));
  INV_X1    g0469(.A(new_n512), .ZN(new_n670));
  NOR4_X1   g0470(.A1(new_n652), .A2(new_n653), .A3(new_n320), .A4(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n663), .B1(new_n519), .B2(new_n522), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n493), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT92), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n668), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n679), .B(new_n609), .C1(new_n666), .C2(new_n667), .ZN(new_n680));
  INV_X1    g0480(.A(new_n665), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n645), .A2(new_n609), .A3(new_n648), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n469), .B1(new_n678), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n463), .A2(new_n464), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n322), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n461), .B2(new_n450), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n413), .A2(new_n414), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n426), .B(new_n428), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n349), .A2(new_n351), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n344), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(G369));
  NAND2_X1  g0493(.A1(new_n296), .A2(new_n227), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n669), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n493), .A2(new_n699), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n657), .A2(new_n673), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n529), .A2(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(KEYINPUT93), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT93), .B1(new_n702), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n699), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n675), .A2(new_n676), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n705), .A2(new_n706), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n575), .B1(new_n560), .B2(new_n708), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n564), .A2(new_n545), .A3(new_n699), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n230), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n225), .A2(new_n721), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n268), .A2(G116), .A3(new_n622), .ZN(new_n723));
  OAI21_X1  g0523(.A(G1), .B1(new_n720), .B2(G41), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  AND4_X1   g0526(.A1(new_n562), .A2(new_n639), .A3(new_n640), .A4(new_n607), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(KEYINPUT30), .A3(new_n654), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n555), .A2(new_n320), .A3(new_n637), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n516), .A2(new_n591), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT30), .B1(new_n727), .B2(new_n654), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT94), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n728), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n509), .A2(new_n515), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n562), .A2(new_n639), .A3(new_n640), .A4(new_n607), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n699), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n650), .A2(new_n530), .A3(new_n575), .A4(new_n708), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n730), .A2(new_n737), .A3(new_n728), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT29), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT95), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n529), .A2(new_n564), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n668), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n619), .A2(new_n524), .ZN(new_n751));
  INV_X1    g0551(.A(new_n667), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n662), .A2(new_n665), .A3(KEYINPUT91), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n673), .A2(new_n669), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n751), .A2(KEYINPUT95), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n665), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n609), .B1(new_n666), .B2(new_n667), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(KEYINPUT26), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n750), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n747), .B1(new_n760), .B2(new_n708), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n527), .A2(new_n528), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT92), .B1(new_n762), .B2(new_n493), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n674), .B(new_n492), .C1(new_n527), .C2(new_n528), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n669), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n754), .A3(new_n751), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n680), .A2(new_n683), .ZN(new_n767));
  AOI211_X1 g0567(.A(KEYINPUT29), .B(new_n699), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n746), .A2(new_n761), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n726), .B1(new_n769), .B2(G1), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT96), .Z(G364));
  AOI21_X1  g0571(.A(new_n226), .B1(G20), .B2(new_n663), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n520), .A2(G20), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(G179), .A3(new_n277), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT100), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n220), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n227), .A2(new_n520), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n780), .A2(new_n277), .A3(G179), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n263), .B1(new_n782), .B2(new_n214), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n320), .A2(new_n277), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n779), .A2(G179), .A3(new_n277), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n786), .A2(new_n207), .B1(new_n201), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n774), .A2(new_n320), .A3(new_n277), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n774), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G179), .A3(new_n277), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n790), .A2(new_n202), .B1(new_n792), .B2(new_n218), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n778), .A2(new_n783), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(KEYINPUT98), .A2(G179), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT98), .B1(G179), .B2(G200), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n520), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n227), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G97), .ZN(new_n801));
  INV_X1    g0601(.A(new_n797), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n791), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT32), .B1(new_n808), .B2(G159), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n808), .A2(KEYINPUT32), .A3(G159), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n794), .B(new_n801), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n387), .B1(new_n782), .B2(new_n552), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n790), .A2(new_n813), .B1(new_n792), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n785), .A2(G326), .ZN(new_n816));
  INV_X1    g0616(.A(G322), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n787), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n812), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n808), .A2(G329), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n800), .A2(G294), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n776), .A2(G283), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n773), .B1(new_n811), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n295), .A2(G20), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n299), .B1(new_n825), .B2(G45), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n721), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n720), .A2(new_n387), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G355), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(G116), .B2(new_n230), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n246), .A2(new_n255), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n720), .A2(new_n263), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n225), .B2(new_n255), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(G13), .A2(G33), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(G20), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n772), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n828), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT97), .Z(new_n843));
  INV_X1    g0643(.A(new_n715), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n824), .B(new_n843), .C1(new_n844), .C2(new_n839), .ZN(new_n845));
  INV_X1    g0645(.A(new_n716), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n828), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n715), .A2(G330), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NAND2_X1  g0651(.A1(new_n773), .A2(new_n838), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n828), .B1(G77), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n777), .A2(new_n214), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n786), .A2(new_n552), .B1(new_n855), .B2(new_n787), .ZN(new_n856));
  INV_X1    g0656(.A(G283), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n790), .A2(new_n857), .B1(new_n792), .B2(new_n477), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n808), .A2(G311), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n263), .B1(new_n781), .B2(G107), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT101), .Z(new_n862));
  NAND4_X1  g0662(.A1(new_n859), .A2(new_n801), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n777), .A2(new_n202), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n387), .B(new_n864), .C1(G50), .C2(new_n781), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n785), .A2(G137), .B1(new_n789), .B2(G150), .ZN(new_n866));
  INV_X1    g0666(.A(new_n787), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(G143), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(new_n399), .C2(new_n792), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT34), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n865), .B(new_n870), .C1(new_n201), .C2(new_n799), .ZN(new_n871));
  INV_X1    g0671(.A(G132), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n807), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n863), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n853), .B1(new_n874), .B2(new_n772), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n309), .A2(new_n699), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n322), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n315), .A2(new_n322), .A3(new_n876), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n875), .B1(new_n879), .B2(new_n838), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n708), .B1(new_n678), .B2(new_n684), .ZN(new_n881));
  INV_X1    g0681(.A(new_n879), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n708), .B(new_n879), .C1(new_n678), .C2(new_n684), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n746), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n828), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n880), .B1(new_n891), .B2(new_n892), .ZN(G384));
  OR2_X1    g0693(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(G116), .A3(new_n228), .A4(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT36), .Z(new_n897));
  OAI211_X1 g0697(.A(new_n225), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n207), .A2(G68), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n299), .B(G13), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n450), .A2(new_n461), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n699), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n383), .A2(new_n410), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(new_n697), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n420), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n905), .A2(new_n425), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n905), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n400), .B1(new_n401), .B2(G20), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n415), .B2(new_n416), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n398), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n911), .B(new_n386), .C1(new_n914), .C2(new_n403), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n408), .B1(new_n390), .B2(new_n396), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n417), .B(new_n280), .C1(new_n916), .C2(KEYINPUT16), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT103), .B1(new_n917), .B2(new_n419), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n370), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n379), .A2(new_n320), .A3(new_n380), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT77), .B1(new_n366), .B2(new_n275), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n697), .B1(new_n923), .B2(new_n422), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n910), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n909), .B1(new_n925), .B2(new_n906), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n915), .A2(new_n918), .A3(new_n697), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n429), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n904), .B(KEYINPUT39), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n908), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n429), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n905), .A2(new_n425), .A3(new_n908), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT37), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n909), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n931), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n928), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n917), .A2(new_n419), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n911), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n917), .A2(KEYINPUT103), .A3(new_n419), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n924), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n906), .B1(new_n948), .B2(new_n905), .ZN(new_n949));
  INV_X1    g0749(.A(new_n909), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n938), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n941), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n904), .B1(new_n953), .B2(KEYINPUT39), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n903), .B1(new_n943), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n907), .B1(new_n426), .B2(new_n428), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n461), .B(new_n699), .C1(new_n686), .C2(new_n450), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n461), .A2(new_n699), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n465), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n322), .A2(new_n699), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n961), .B1(new_n885), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n956), .B1(new_n964), .B2(new_n953), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n955), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n469), .B1(new_n761), .B2(new_n768), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n692), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(KEYINPUT31), .B(new_n699), .C1(new_n733), .C2(new_n738), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n741), .A2(new_n742), .A3(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n957), .A2(new_n959), .B1(new_n878), .B2(new_n877), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n929), .C2(new_n930), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n971), .A2(new_n972), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT40), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n939), .B2(new_n941), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n973), .A2(new_n975), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n469), .A3(new_n971), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(G330), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n979), .B1(new_n469), .B2(new_n971), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n969), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n299), .B2(new_n825), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n969), .A2(new_n983), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n901), .B1(new_n985), .B2(new_n986), .ZN(G367));
  INV_X1    g0787(.A(new_n707), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n660), .B1(new_n606), .B2(new_n708), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n609), .A2(new_n699), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n615), .A2(new_n618), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n610), .B1(new_n993), .B2(new_n673), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n992), .A2(KEYINPUT42), .B1(new_n708), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n991), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n707), .A2(KEYINPUT42), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n665), .A2(new_n629), .A3(new_n708), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n629), .A2(new_n708), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n754), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n717), .A2(new_n991), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n995), .A2(new_n1002), .A3(new_n1001), .A4(new_n997), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n721), .B(KEYINPUT41), .Z(new_n1012));
  NAND3_X1  g0812(.A1(new_n707), .A2(new_n709), .A3(new_n991), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1013), .B(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT44), .B1(new_n710), .B2(new_n996), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT44), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1018), .B(new_n991), .C1(new_n707), .C2(new_n709), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n717), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1013), .B(new_n1014), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1022), .B(new_n718), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n746), .A2(new_n761), .A3(new_n768), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n705), .A2(new_n706), .A3(new_n700), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n716), .B1(new_n988), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1025), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1027), .A2(new_n707), .A3(new_n846), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1021), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1012), .B1(new_n1031), .B2(new_n769), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1011), .B1(new_n1032), .B2(new_n827), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n242), .A2(new_n833), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1034), .B(new_n840), .C1(new_n230), .C2(new_n287), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n792), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1036), .A2(G50), .B1(new_n789), .B2(G159), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1038), .A2(KEYINPUT108), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(KEYINPUT108), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n781), .A2(G58), .B1(new_n785), .B2(G143), .ZN(new_n1041));
  INV_X1    g0841(.A(G150), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n787), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1039), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n808), .A2(G137), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n387), .B1(new_n775), .B2(G77), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT109), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n800), .A2(G68), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT46), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n782), .B2(new_n477), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n855), .C2(new_n790), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT107), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n387), .B1(new_n792), .B2(new_n857), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n775), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1056), .A2(new_n593), .B1(new_n552), .B2(new_n787), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G311), .C2(new_n785), .ZN(new_n1058));
  INV_X1    g0858(.A(G317), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n807), .C1(new_n269), .C2(new_n799), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT47), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n828), .B(new_n1035), .C1(new_n1062), .C2(new_n773), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT110), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1001), .A2(new_n839), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1033), .A2(new_n1066), .ZN(G387));
  OR2_X1    g0867(.A1(new_n239), .A2(new_n255), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1068), .A2(new_n833), .B1(new_n723), .B2(new_n829), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n336), .B2(new_n207), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n255), .B1(new_n202), .B2(new_n218), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n723), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1069), .A2(new_n1074), .B1(G107), .B2(new_n230), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n890), .B1(new_n1075), .B2(new_n840), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n799), .A2(new_n287), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n786), .A2(new_n399), .B1(new_n207), .B2(new_n787), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n387), .B(new_n1078), .C1(G77), .C2(new_n781), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1036), .A2(G68), .B1(new_n789), .B2(new_n336), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT111), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(new_n593), .C2(new_n777), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1077), .B(new_n1082), .C1(G150), .C2(new_n808), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n785), .A2(G322), .B1(new_n789), .B2(G311), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n552), .B2(new_n792), .C1(new_n1059), .C2(new_n787), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT112), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n800), .A2(G283), .B1(G294), .B2(new_n781), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n808), .A2(G326), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n387), .B1(new_n1056), .B2(new_n477), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1083), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1076), .B1(new_n1098), .B2(new_n773), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n712), .B2(new_n839), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1029), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n827), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n769), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n721), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(G393));
  NAND2_X1  g0905(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1030), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n721), .A3(new_n1031), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1021), .A2(new_n1023), .A3(new_n827), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n996), .A2(new_n839), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n263), .B1(new_n792), .B2(new_n289), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n782), .A2(new_n202), .B1(new_n790), .B2(new_n207), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n854), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n808), .A2(G143), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n800), .A2(G77), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n786), .A2(new_n1042), .B1(new_n399), .B2(new_n787), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT51), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n263), .B(new_n778), .C1(G283), .C2(new_n781), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n786), .A2(new_n1059), .B1(new_n814), .B2(new_n787), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT52), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1120), .B(new_n1122), .C1(new_n817), .C2(new_n807), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1036), .A2(G294), .B1(new_n789), .B2(G303), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n799), .B2(new_n477), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT113), .Z(new_n1126));
  OAI21_X1  g0926(.A(new_n1119), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n772), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n840), .B1(new_n593), .B2(new_n230), .C1(new_n249), .C2(new_n834), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1111), .A2(new_n828), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1110), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1109), .A2(new_n1131), .ZN(G390));
  OAI21_X1  g0932(.A(KEYINPUT39), .B1(new_n929), .B2(new_n930), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT104), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n942), .A3(new_n931), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n885), .A2(new_n963), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n903), .B1(new_n1136), .B2(new_n960), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n760), .A2(new_n708), .A3(new_n879), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n961), .B1(new_n1138), .B2(new_n963), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n939), .A2(new_n941), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n902), .B2(new_n699), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1135), .A2(new_n1137), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n971), .A2(G330), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1143), .A2(new_n882), .A3(new_n961), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1143), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n469), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n967), .A2(new_n692), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n960), .B1(new_n746), .B2(new_n879), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1136), .B1(new_n1149), .B2(new_n1144), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n746), .A2(new_n879), .A3(new_n960), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n961), .B1(new_n1143), .B2(new_n882), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1151), .A2(new_n963), .A3(new_n1152), .A4(new_n1138), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1148), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1151), .B1(new_n1139), .B2(new_n1141), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1145), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(KEYINPUT114), .A3(new_n721), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1145), .A2(new_n1155), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT114), .B1(new_n1156), .B2(new_n721), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1145), .A2(new_n827), .A3(new_n1155), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT116), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n828), .B1(new_n336), .B2(new_n852), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n807), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n792), .A2(new_n1168), .B1(new_n787), .B2(new_n872), .ZN(new_n1169));
  INV_X1    g0969(.A(G128), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n786), .A2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G137), .C2(new_n789), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT53), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n782), .B2(new_n1042), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n781), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n263), .B1(new_n1056), .B2(new_n207), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT115), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1174), .A2(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n800), .A2(G159), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1172), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n864), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n263), .B1(new_n781), .B2(G87), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n786), .A2(new_n857), .B1(new_n593), .B2(new_n792), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n790), .A2(new_n269), .B1(new_n477), .B2(new_n787), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1182), .A2(new_n1116), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n807), .A2(new_n855), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1167), .A2(new_n1181), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1165), .B1(new_n1189), .B2(new_n772), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1135), .B2(new_n838), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1163), .A2(new_n1164), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1164), .B1(new_n1163), .B2(new_n1191), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1161), .A2(new_n1162), .B1(new_n1192), .B2(new_n1193), .ZN(G378));
  INV_X1    g0994(.A(new_n1148), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1156), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n343), .A2(new_n697), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT119), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n352), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n352), .A2(new_n1199), .ZN(new_n1201));
  XOR2_X1   g1001(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR3_X1    g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n979), .B2(G330), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n973), .A2(new_n975), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n978), .A2(new_n971), .A3(new_n972), .ZN(new_n1209));
  AND4_X1   g1009(.A1(G330), .A2(new_n1208), .A3(new_n1209), .A4(new_n1206), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n966), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(G330), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1206), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1208), .A2(new_n1209), .A3(G330), .A4(new_n1206), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(new_n955), .A3(new_n965), .A4(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1211), .A2(KEYINPUT57), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1196), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1195), .B2(new_n1156), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n721), .C1(new_n1220), .C2(KEYINPUT57), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1211), .A2(new_n1216), .A3(new_n827), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n828), .B1(G50), .B2(new_n852), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n254), .B(new_n387), .C1(new_n782), .C2(new_n218), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT117), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n201), .B2(new_n1056), .C1(new_n857), .C2(new_n807), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT118), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n867), .A2(G107), .B1(G97), .B2(new_n789), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n287), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1036), .A2(new_n1229), .B1(G116), .B2(new_n785), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1048), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT58), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G33), .A2(G41), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G50), .B(new_n1235), .C1(new_n387), .C2(new_n254), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n782), .A2(new_n1168), .B1(new_n786), .B2(new_n1166), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G137), .B2(new_n1036), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n867), .A2(G128), .B1(G132), .B2(new_n789), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n1042), .C2(new_n799), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1241));
  INV_X1    g1041(.A(G124), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1235), .B1(new_n399), .B2(new_n1056), .C1(new_n807), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1240), .B2(KEYINPUT59), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1236), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1233), .A2(new_n1234), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1223), .B1(new_n1246), .B2(new_n772), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n838), .B2(new_n1213), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1222), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1221), .A2(new_n1250), .ZN(G375));
  NAND2_X1  g1051(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n961), .A2(new_n837), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n828), .B1(G68), .B2(new_n852), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n387), .B1(new_n775), .B2(G58), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT120), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n790), .A2(new_n1168), .B1(new_n792), .B2(new_n1042), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n867), .A2(G137), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n782), .A2(new_n399), .B1(new_n786), .B2(new_n872), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n207), .B2(new_n799), .C1(new_n1170), .C2(new_n807), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n807), .A2(new_n552), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n782), .A2(new_n593), .B1(new_n269), .B2(new_n792), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n786), .A2(new_n855), .B1(new_n857), .B2(new_n787), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n387), .B1(new_n790), .B2(new_n477), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n218), .B2(new_n777), .C1(new_n287), .C2(new_n799), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1254), .B1(new_n1268), .B2(new_n772), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1252), .A2(new_n827), .B1(new_n1253), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1012), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1159), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1252), .A2(new_n1195), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1270), .B1(new_n1272), .B2(new_n1273), .ZN(G381));
  OAI211_X1 g1074(.A(new_n1102), .B(new_n850), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1275), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G387), .A2(new_n1276), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n698), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  NAND2_X1  g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1275), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1284), .A2(new_n1109), .A3(new_n1131), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1109), .B2(new_n1131), .ZN(new_n1286));
  OAI21_X1  g1086(.A(G387), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G390), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1284), .A2(new_n1109), .A3(new_n1131), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1289), .A2(new_n1033), .A3(new_n1066), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G378), .A2(new_n1221), .A3(new_n1250), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT121), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1249), .A2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1196), .A2(new_n1271), .A3(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1222), .A2(KEYINPUT121), .A3(new_n1248), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1162), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1193), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1163), .A2(new_n1164), .A3(new_n1191), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1299), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1293), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT122), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT123), .ZN(new_n1308));
  OR2_X1    g1108(.A1(G384), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1270), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G384), .A2(new_n1308), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1273), .B1(KEYINPUT60), .B2(new_n1159), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1150), .A2(new_n1148), .A3(new_n1153), .A4(KEYINPUT60), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n721), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1311), .B(new_n1312), .C1(new_n1313), .C2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1312), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(new_n1310), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT122), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1293), .A2(new_n1305), .A3(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1307), .A2(new_n1279), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1280), .B1(new_n1293), .B2(new_n1305), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1320), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(new_n1324), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1323), .A2(new_n1324), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1280), .A2(G2897), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT124), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1280), .A2(KEYINPUT124), .A3(G2897), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1320), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1316), .A2(new_n1331), .A3(new_n1319), .A4(new_n1330), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1329), .B1(new_n1337), .B2(new_n1325), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1292), .B1(new_n1328), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1323), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1307), .A2(new_n1279), .A3(new_n1322), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1336), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1340), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1306), .A2(new_n1279), .A3(new_n1344), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1287), .A2(new_n1291), .A3(new_n1329), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  AND4_X1   g1148(.A1(KEYINPUT125), .A2(new_n1341), .A3(new_n1343), .A4(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1347), .B1(new_n1342), .B2(new_n1336), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT125), .B1(new_n1350), .B2(new_n1341), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1339), .B1(new_n1349), .B2(new_n1351), .ZN(G405));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1278), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1326), .A2(new_n1353), .A3(new_n1293), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1354), .B(KEYINPUT127), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT126), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1293), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1356), .B1(new_n1357), .B2(new_n1320), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1357), .A2(new_n1356), .A3(new_n1320), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1355), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1292), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1292), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1355), .B(new_n1362), .C1(new_n1358), .C2(new_n1359), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1361), .A2(new_n1363), .ZN(G402));
endmodule


