//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT74), .B(G211gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT22), .B1(new_n207), .B2(G218gat), .ZN(new_n208));
  XOR2_X1   g007(.A(G197gat), .B(G204gat), .Z(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT74), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G211gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n214), .A3(G218gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT22), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n209), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n205), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT23), .B(new_n221), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n224), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT23), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n232), .A3(new_n233), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n234), .A2(new_n246), .A3(new_n235), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n245), .A2(new_n239), .A3(new_n240), .A4(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n248), .A2(new_n232), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n237), .B2(KEYINPUT69), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n256), .ZN(new_n258));
  NAND3_X1  g057(.A1(KEYINPUT68), .A2(KEYINPUT27), .A3(G183gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n238), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n227), .A2(new_n265), .A3(KEYINPUT26), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT26), .B1(new_n227), .B2(new_n265), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n233), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n261), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n252), .A2(new_n253), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n244), .A2(new_n271), .A3(new_n251), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n244), .B2(new_n251), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n253), .A2(KEYINPUT29), .ZN(new_n275));
  AOI211_X1 g074(.A(new_n220), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n220), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n253), .B(new_n269), .C1(new_n272), .C2(new_n273), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n252), .A2(new_n269), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n276), .A2(KEYINPUT75), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(new_n275), .ZN(new_n284));
  INV_X1    g083(.A(new_n270), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n277), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n220), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n283), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n204), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n204), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n281), .B1(new_n277), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT30), .A3(new_n291), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT39), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(G148gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n310), .B2(KEYINPUT2), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(G141gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n313), .A2(new_n305), .B1(KEYINPUT76), .B2(KEYINPUT2), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT77), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G155gat), .B2(G162gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n315), .A2(new_n317), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G127gat), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G113gat), .B(G120gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(KEYINPUT1), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n329), .A2(new_n337), .A3(KEYINPUT79), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT79), .B1(new_n329), .B2(new_n337), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n322), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND4_X1   g139(.A1(new_n319), .A2(new_n315), .A3(new_n317), .A4(new_n320), .ZN(new_n341));
  INV_X1    g140(.A(new_n314), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n342), .B1(new_n311), .B2(new_n306), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n329), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n299), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n312), .B(new_n349), .C1(new_n314), .C2(new_n321), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT80), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n341), .A2(new_n342), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n349), .A4(new_n312), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n337), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n329), .A2(new_n337), .A3(KEYINPUT79), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(new_n322), .B2(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n344), .A3(new_n362), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n355), .A2(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n348), .B1(new_n347), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT85), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(G57gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  INV_X1    g168(.A(G85gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n368), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n362), .B1(new_n343), .B2(new_n344), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n322), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n347), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n299), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n365), .A2(new_n372), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT40), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n378), .A3(KEYINPUT40), .A4(new_n372), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n346), .B2(new_n347), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n340), .A2(new_n345), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT83), .A3(new_n377), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(KEYINPUT81), .B(KEYINPUT4), .C1(new_n322), .C2(new_n356), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n347), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n375), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT82), .B1(new_n394), .B2(new_n373), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n361), .A2(new_n393), .A3(new_n363), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n377), .B1(new_n374), .B2(KEYINPUT81), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n373), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n389), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n376), .A2(KEYINPUT5), .A3(new_n377), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n372), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n383), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n210), .B2(new_n219), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n322), .B1(new_n407), .B2(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n351), .B2(new_n354), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n220), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n409), .B2(new_n220), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n413), .ZN(new_n415));
  OAI221_X1 g214(.A(new_n408), .B1(new_n411), .B2(new_n415), .C1(new_n409), .C2(new_n220), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n406), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(new_n406), .A3(new_n416), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT31), .B(G50gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n422), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n418), .B(new_n424), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n419), .A2(new_n423), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n419), .B2(new_n425), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n417), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n298), .A2(new_n405), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT37), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT75), .B1(new_n276), .B2(new_n281), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n286), .A2(new_n288), .A3(new_n283), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n286), .A2(new_n288), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n204), .B1(new_n437), .B2(KEYINPUT37), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT38), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n372), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT83), .B1(new_n387), .B2(new_n377), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n385), .B(new_n347), .C1(new_n340), .C2(new_n345), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT5), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n398), .A2(new_n399), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n394), .A2(KEYINPUT82), .A3(new_n373), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT6), .B(new_n440), .C1(new_n446), .C2(new_n402), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n440), .B1(new_n446), .B2(new_n402), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n401), .A2(new_n372), .A3(new_n403), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n292), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n291), .A2(KEYINPUT38), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n296), .B2(new_n433), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n433), .B1(new_n287), .B2(new_n277), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n295), .A2(new_n220), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n439), .A2(new_n447), .A3(new_n451), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n432), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n447), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n297), .A2(new_n294), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n291), .B1(new_n434), .B2(new_n435), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n428), .A2(new_n431), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G227gat), .ZN(new_n469));
  INV_X1    g268(.A(G233gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n244), .A2(new_n271), .A3(new_n251), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n344), .B1(new_n474), .B2(new_n269), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n344), .B(new_n269), .C1(new_n272), .C2(new_n273), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G15gat), .B(G43gat), .Z(new_n482));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n274), .A2(new_n356), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n476), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n488), .B2(new_n471), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n490), .A2(KEYINPUT33), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT72), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n471), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n487), .B2(new_n476), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497));
  NOR4_X1   g296(.A1(new_n496), .A2(new_n497), .A3(new_n486), .A4(new_n492), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n485), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n487), .A2(new_n495), .A3(new_n476), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n502), .B(new_n485), .C1(new_n494), .C2(new_n498), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(KEYINPUT36), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT36), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n460), .B(new_n468), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n466), .A3(new_n505), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n504), .A2(new_n466), .A3(KEYINPUT89), .A4(new_n505), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n461), .A2(new_n464), .A3(KEYINPUT35), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n509), .B2(new_n465), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n508), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI221_X1 g324(.A(new_n521), .B1(new_n522), .B2(new_n518), .C1(G1gat), .C2(new_n519), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT97), .ZN(new_n529));
  XOR2_X1   g328(.A(G57gat), .B(G64gat), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G71gat), .B(G78gat), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n532), .ZN(new_n534));
  NAND3_X1  g333(.A1(KEYINPUT98), .A2(G57gat), .A3(G64gat), .ZN(new_n535));
  AND2_X1   g334(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(G64gat), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n529), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n527), .B1(new_n539), .B2(KEYINPUT21), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n546));
  XNOR2_X1  g345(.A(G183gat), .B(G211gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT99), .ZN(new_n549));
  OR3_X1    g348(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n544), .B2(new_n545), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n552));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n550), .B2(new_n551), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n370), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n370), .B2(new_n559), .ZN(new_n562));
  NAND3_X1  g361(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G99gat), .B(G106gat), .Z(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT102), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(KEYINPUT102), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT14), .ZN(new_n573));
  NOR2_X1   g372(.A1(G29gat), .A2(G36gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(KEYINPUT90), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(KEYINPUT90), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT15), .ZN(new_n578));
  XOR2_X1   g377(.A(G43gat), .B(G50gat), .Z(new_n579));
  XOR2_X1   g378(.A(KEYINPUT91), .B(G29gat), .Z(new_n580));
  AOI22_X1  g379(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(G36gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n579), .A2(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n577), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n584), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT93), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT17), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n584), .B2(new_n586), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n597), .A2(KEYINPUT103), .A3(new_n572), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT103), .B1(new_n597), .B2(new_n572), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n589), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT101), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n601), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n607), .B(new_n589), .C1(new_n598), .C2(new_n599), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n606), .B1(new_n602), .B2(new_n608), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n557), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  INV_X1    g413(.A(new_n527), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n591), .B2(new_n595), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n584), .A2(new_n586), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n527), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n619), .B(new_n615), .C1(new_n591), .C2(new_n595), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT18), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n614), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G113gat), .B(G141gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G197gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT11), .B(G169gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  NOR2_X1   g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n617), .B(new_n527), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n623), .B(KEYINPUT13), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n626), .A2(new_n627), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n621), .A2(KEYINPUT18), .A3(new_n624), .A4(new_n625), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n638), .B(new_n639), .C1(new_n628), .C2(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n533), .A2(new_n538), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n568), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n533), .A2(new_n538), .A3(new_n566), .A4(new_n567), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n570), .A2(new_n539), .A3(KEYINPUT10), .A4(new_n571), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n648), .B2(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n654), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n656), .A2(KEYINPUT105), .A3(new_n654), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT106), .B1(new_n655), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n649), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n654), .B1(new_n667), .B2(KEYINPUT104), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n664), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n654), .B1(new_n648), .B2(new_n649), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n662), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n643), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n613), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n517), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT107), .ZN(new_n683));
  INV_X1    g482(.A(new_n461), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n298), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n688), .A2(KEYINPUT108), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT108), .B1(new_n688), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n518), .B1(new_n683), .B2(new_n298), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n693), .B2(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n504), .A2(new_n505), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(G15gat), .B1(new_n683), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n506), .A2(new_n507), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n698), .B1(new_n683), .B2(new_n701), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n467), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(new_n611), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n609), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n517), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n680), .A2(new_n557), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n461), .A3(new_n580), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT45), .Z(new_n712));
  AOI21_X1  g511(.A(new_n298), .B1(new_n447), .B2(new_n451), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT109), .B1(new_n713), .B2(new_n466), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n465), .A2(new_n715), .A3(new_n467), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n460), .B1(new_n506), .B2(new_n507), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n516), .B(new_n514), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n719), .B2(new_n707), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n517), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT110), .B1(new_n722), .B2(new_n709), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  INV_X1    g524(.A(new_n709), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n720), .A2(new_n721), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n461), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n580), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n712), .B1(new_n729), .B2(new_n730), .ZN(G1328gat));
  NOR3_X1   g530(.A1(new_n710), .A2(G36gat), .A3(new_n464), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT46), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n464), .B1(new_n724), .B2(new_n728), .ZN(new_n734));
  INV_X1    g533(.A(G36gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n721), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n707), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n726), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n700), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n710), .A2(G43gat), .A3(new_n696), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n700), .B1(new_n723), .B2(new_n727), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g550(.A1(new_n742), .A2(new_n467), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G50gat), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n710), .A2(G50gat), .A3(new_n466), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n467), .B1(new_n723), .B2(new_n727), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n754), .B1(new_n758), .B2(G50gat), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n760));
  OAI21_X1  g559(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(G1331gat));
  NOR3_X1   g560(.A1(new_n613), .A2(new_n643), .A3(new_n679), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n719), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(KEYINPUT112), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n684), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  OAI22_X1  g568(.A1(new_n766), .A2(new_n464), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT49), .B(G64gat), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n764), .A2(new_n298), .A3(new_n765), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n771), .B1(new_n770), .B2(new_n773), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(G1333gat));
  NAND4_X1  g576(.A1(new_n764), .A2(G71gat), .A3(new_n700), .A4(new_n765), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n766), .A2(new_n696), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(G71gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n778), .B(new_n782), .C1(new_n779), .C2(G71gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n467), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n557), .A2(new_n643), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n719), .A2(new_n707), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n679), .A2(new_n461), .A3(G85gat), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT116), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n787), .A2(new_n678), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT114), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n722), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n684), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n795), .B1(new_n370), .B2(new_n799), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n722), .A2(new_n298), .A3(new_n797), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n801), .A2(G92gat), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n790), .A2(new_n559), .A3(new_n298), .A4(new_n678), .ZN(new_n803));
  OR2_X1    g602(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n802), .B2(new_n803), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(G1337gat));
  NOR3_X1   g606(.A1(new_n696), .A2(G99gat), .A3(new_n679), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n798), .A2(new_n700), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G99gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1338gat));
  NOR2_X1   g611(.A1(new_n466), .A2(G106gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n678), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n722), .A2(new_n467), .A3(new_n797), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g617(.A1(new_n511), .A2(new_n512), .ZN(new_n819));
  INV_X1    g618(.A(new_n557), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n670), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n676), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n662), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n822), .B1(new_n668), .B2(new_n669), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT55), .B1(new_n831), .B2(new_n827), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n830), .A2(new_n832), .B1(new_n666), .B2(new_n673), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n643), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n632), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n624), .B1(new_n621), .B2(new_n625), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n635), .A2(new_n637), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n638), .A2(new_n633), .A3(new_n639), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n678), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n707), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n833), .B1(new_n610), .B2(new_n611), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n841), .A3(new_n840), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n820), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n643), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n679), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n613), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n819), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n461), .A2(new_n298), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n332), .A3(new_n643), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n847), .A2(new_n851), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n466), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT119), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(new_n697), .A3(new_n643), .A4(new_n853), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(KEYINPUT120), .A3(G113gat), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT120), .B1(new_n859), .B2(G113gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n855), .B1(new_n860), .B2(new_n861), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n697), .A3(new_n853), .ZN(new_n863));
  OAI21_X1  g662(.A(G120gat), .B1(new_n863), .B2(new_n679), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n854), .A2(new_n330), .A3(new_n678), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  NOR3_X1   g665(.A1(new_n863), .A2(new_n325), .A3(new_n820), .ZN(new_n867));
  AOI21_X1  g666(.A(G127gat), .B1(new_n854), .B2(new_n557), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1342gat));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n323), .A3(new_n707), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT56), .Z(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n863), .B2(new_n612), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1343gat));
  AND2_X1   g672(.A1(new_n699), .A2(new_n853), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n466), .B1(new_n847), .B2(new_n851), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n829), .B1(new_n824), .B2(new_n828), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n674), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n642), .B2(new_n641), .ZN(new_n880));
  AND4_X1   g679(.A1(new_n678), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n612), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n845), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n707), .A2(new_n883), .A3(new_n833), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n557), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT57), .B(new_n467), .C1(new_n885), .C2(new_n850), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n856), .B2(new_n467), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n874), .B(new_n876), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890), .B2(new_n848), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n874), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n301), .A3(new_n643), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n897), .A3(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n891), .B(new_n896), .C1(new_n892), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n303), .A3(new_n678), .ZN(new_n902));
  INV_X1    g701(.A(new_n890), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n303), .C1(new_n903), .C2(new_n678), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n844), .A2(KEYINPUT123), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n845), .B1(new_n844), .B2(KEYINPUT123), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n843), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n851), .B1(new_n908), .B2(new_n557), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n467), .ZN(new_n910));
  INV_X1    g709(.A(new_n886), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n678), .B(new_n874), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n905), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n902), .B1(new_n904), .B2(new_n913), .ZN(G1345gat));
  AOI21_X1  g713(.A(G155gat), .B1(new_n895), .B2(new_n557), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n820), .A2(new_n308), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n903), .B2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n890), .B2(new_n612), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n309), .A3(new_n707), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n684), .A2(new_n464), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n857), .A2(KEYINPUT119), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n856), .B2(new_n466), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n697), .B(new_n921), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n848), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n852), .A2(new_n921), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n221), .A3(new_n643), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1348gat));
  OR3_X1    g728(.A1(new_n679), .A2(new_n223), .A3(new_n225), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n927), .A2(new_n678), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n925), .A2(new_n930), .B1(new_n931), .B2(G176gat), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n925), .B2(new_n820), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n557), .A2(new_n262), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT125), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n238), .A3(new_n707), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  NAND4_X1  g746(.A1(new_n858), .A2(new_n697), .A3(new_n707), .A4(new_n921), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n948), .B2(G190gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  AND2_X1   g751(.A1(new_n699), .A2(new_n921), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n875), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  XOR2_X1   g754(.A(KEYINPUT127), .B(G197gat), .Z(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n643), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n910), .A2(new_n911), .ZN(new_n958));
  INV_X1    g757(.A(new_n953), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n958), .A2(new_n848), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n960), .B2(new_n956), .ZN(G1352gat));
  NOR3_X1   g760(.A1(new_n954), .A2(G204gat), .A3(new_n679), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n958), .A2(new_n679), .A3(new_n959), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G1353gat));
  OR3_X1    g765(.A1(new_n954), .A2(new_n207), .A3(new_n820), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n557), .B(new_n953), .C1(new_n910), .C2(new_n911), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  AOI21_X1  g770(.A(G218gat), .B1(new_n955), .B2(new_n707), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n958), .A2(new_n959), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n707), .A2(G218gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1355gat));
endmodule


