//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207));
  OAI21_X1  g006(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n208), .B(new_n209), .Z(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n210), .B1(new_n219), .B2(KEYINPUT66), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(KEYINPUT66), .B2(new_n219), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT24), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(KEYINPUT24), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT68), .B(G190gat), .Z(new_n230));
  OAI211_X1 g029(.A(new_n228), .B(new_n229), .C1(G183gat), .C2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n218), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n232), .A4(new_n212), .ZN(new_n233));
  INV_X1    g032(.A(new_n230), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT28), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT27), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(KEYINPUT69), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n225), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(KEYINPUT70), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(KEYINPUT70), .ZN(new_n244));
  AOI211_X1 g043(.A(new_n230), .B(new_n238), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n236), .B1(new_n245), .B2(KEYINPUT28), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n225), .A2(new_n226), .ZN(new_n247));
  INV_X1    g046(.A(G169gat), .ZN(new_n248));
  INV_X1    g047(.A(G176gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n250), .A2(KEYINPUT26), .A3(new_n211), .ZN(new_n251));
  AOI211_X1 g050(.A(new_n247), .B(new_n251), .C1(KEYINPUT26), .C2(new_n211), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n223), .A2(new_n233), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n207), .B1(new_n253), .B2(KEYINPUT29), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n223), .A2(new_n233), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n246), .A2(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n207), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260));
  INV_X1    g059(.A(G211gat), .ZN(new_n261));
  INV_X1    g060(.A(G218gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(KEYINPUT22), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G211gat), .B(G218gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(KEYINPUT73), .A3(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n259), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n273));
  INV_X1    g072(.A(new_n256), .ZN(new_n274));
  INV_X1    g073(.A(new_n233), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n221), .B2(new_n222), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n207), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n270), .B1(new_n278), .B2(new_n259), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n206), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n258), .B1(new_n257), .B2(new_n273), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n207), .B1(new_n255), .B2(new_n256), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n269), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n271), .A3(new_n205), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n284), .A3(KEYINPUT30), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n283), .A2(new_n286), .A3(new_n271), .A4(new_n205), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G1gat), .B(G29gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT0), .ZN(new_n290));
  XNOR2_X1  g089(.A(G57gat), .B(G85gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n290), .B(new_n291), .Z(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G120gat), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n293), .B2(new_n294), .ZN(new_n296));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT71), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G120gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n295), .B(new_n297), .C1(new_n301), .C2(new_n293), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G155gat), .B(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(KEYINPUT2), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n304), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(G162gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(G155gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n307), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT4), .B1(new_n303), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  INV_X1    g114(.A(new_n313), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n315), .A3(new_n316), .A4(new_n302), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G225gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n313), .B(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n321), .B(new_n303), .C1(new_n323), .C2(new_n320), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n303), .A2(new_n313), .ZN(new_n326));
  INV_X1    g125(.A(new_n323), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n303), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n325), .B(KEYINPUT5), .C1(new_n319), .C2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n318), .A2(new_n324), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n319), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n292), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT6), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n329), .A2(new_n332), .A3(new_n292), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(KEYINPUT77), .A3(new_n337), .ZN(new_n341));
  INV_X1    g140(.A(new_n333), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n335), .B1(new_n343), .B2(KEYINPUT78), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n340), .A2(new_n345), .A3(new_n341), .A4(new_n342), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n288), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n255), .A2(new_n303), .A3(new_n256), .ZN(new_n348));
  INV_X1    g147(.A(new_n303), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n274), .B2(new_n276), .ZN(new_n350));
  INV_X1    g149(.A(G227gat), .ZN(new_n351));
  INV_X1    g150(.A(G233gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G15gat), .B(G43gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n348), .A2(new_n350), .ZN(new_n361));
  INV_X1    g160(.A(new_n353), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT34), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT34), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n360), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n354), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n359), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n354), .B2(new_n355), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n365), .B1(new_n361), .B2(new_n362), .ZN(new_n373));
  AOI211_X1 g172(.A(KEYINPUT34), .B(new_n353), .C1(new_n348), .C2(new_n350), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n367), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n367), .B2(new_n375), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n321), .A2(new_n273), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n269), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT79), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n266), .A2(new_n273), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n313), .B1(new_n381), .B2(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n269), .A2(new_n385), .A3(new_n378), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n380), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n320), .B1(new_n269), .B2(KEYINPUT29), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n388), .A2(new_n327), .B1(new_n269), .B2(new_n378), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n383), .ZN(new_n390));
  INV_X1    g189(.A(G22gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G78gat), .B(G106gat), .Z(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT31), .B(G50gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT80), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n387), .B(G22gat), .C1(new_n389), .C2(new_n383), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n395), .A2(KEYINPUT80), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n392), .B2(new_n397), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n376), .A2(new_n377), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n202), .B1(new_n347), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n367), .A2(new_n375), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n401), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n367), .A2(new_n370), .A3(new_n375), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n285), .A2(new_n287), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n342), .A2(new_n337), .A3(new_n336), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT35), .B1(new_n411), .B2(new_n334), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n205), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n282), .B1(new_n207), .B2(new_n277), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n271), .B1(new_n417), .B2(new_n270), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n206), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n283), .B2(new_n271), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT38), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n284), .B(new_n334), .C1(new_n338), .C2(new_n333), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT38), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n254), .A2(new_n259), .A3(new_n269), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(KEYINPUT37), .C1(new_n417), .C2(new_n269), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n205), .B1(new_n283), .B2(new_n271), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n424), .B(new_n426), .C1(new_n427), .C2(new_n416), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT39), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n328), .B2(new_n319), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n319), .B2(new_n330), .ZN(new_n432));
  INV_X1    g231(.A(new_n292), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n319), .B1(new_n318), .B2(new_n324), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n430), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n333), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT40), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n287), .A4(new_n285), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n429), .A2(new_n407), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT36), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n376), .B2(new_n377), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n406), .A2(KEYINPUT36), .A3(new_n408), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n346), .A3(new_n334), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n407), .B1(new_n450), .B2(new_n410), .ZN(new_n451));
  OAI22_X1  g250(.A1(new_n403), .A2(new_n414), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G229gat), .A2(G233gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n453), .B(KEYINPUT13), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G50gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G43gat), .ZN(new_n457));
  INV_X1    g256(.A(G43gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G50gat), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT15), .ZN(new_n460));
  INV_X1    g259(.A(G36gat), .ZN(new_n461));
  INV_X1    g260(.A(G29gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G29gat), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n461), .A3(KEYINPUT14), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(G29gat), .B2(G36gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n460), .B(KEYINPUT85), .C1(new_n466), .C2(new_n470), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT84), .B(G29gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n469), .B(new_n467), .C1(new_n475), .C2(new_n461), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT15), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n459), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(KEYINPUT86), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT86), .A3(new_n477), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n473), .A2(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n391), .A2(G15gat), .ZN(new_n483));
  INV_X1    g282(.A(G15gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G22gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G1gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(KEYINPUT16), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n483), .A2(new_n485), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n483), .A2(new_n485), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT89), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(new_n489), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n488), .A2(new_n496), .A3(new_n494), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n493), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT93), .B1(new_n482), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n474), .ZN(new_n502));
  INV_X1    g301(.A(new_n479), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n466), .A2(new_n470), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n481), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n493), .A2(new_n495), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n498), .A2(new_n499), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n502), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n500), .A3(KEYINPUT93), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n455), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512));
  INV_X1    g311(.A(new_n474), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT85), .B1(new_n476), .B2(new_n460), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n505), .B(KEYINPUT17), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n500), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n482), .B2(KEYINPUT17), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT87), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n512), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(KEYINPUT17), .B2(new_n482), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n517), .B(KEYINPUT17), .C1(new_n502), .C2(new_n505), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT87), .B1(new_n519), .B2(new_n520), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n524), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n511), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n524), .A2(new_n453), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n522), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n530), .A2(KEYINPUT90), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G169gat), .B(G197gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT12), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n540), .A3(new_n547), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n541), .A2(KEYINPUT94), .A3(new_n550), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n452), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT101), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n518), .A2(new_n521), .ZN(new_n564));
  XOR2_X1   g363(.A(G99gat), .B(G106gat), .Z(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI211_X1 g370(.A(KEYINPUT102), .B(new_n565), .C1(new_n567), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n565), .A2(KEYINPUT102), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n565), .A2(KEYINPUT102), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n575), .A2(new_n567), .A3(new_n576), .A4(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(new_n482), .B2(KEYINPUT17), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT103), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT104), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n578), .A2(new_n519), .B1(KEYINPUT41), .B2(new_n560), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n580), .A2(new_n581), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT103), .B1(new_n564), .B2(new_n579), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n584), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n563), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(new_n591), .A3(new_n563), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n599));
  OR2_X1    g398(.A1(G57gat), .A2(G64gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G57gat), .A2(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n602), .B2(KEYINPUT96), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n596), .A2(new_n597), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n598), .A2(new_n603), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n602), .A2(new_n599), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n596), .A2(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n596), .A2(KEYINPUT95), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n500), .B1(new_n619), .B2(new_n612), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n622));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT99), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT98), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n624), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n621), .B2(new_n622), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n618), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n618), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n576), .A2(new_n567), .A3(new_n571), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n574), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n611), .B(new_n607), .C1(new_n636), .C2(new_n572), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n612), .A2(new_n573), .A3(new_n577), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n578), .A2(new_n613), .A3(KEYINPUT10), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n638), .ZN(new_n645));
  INV_X1    g444(.A(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n644), .A2(new_n647), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n595), .A2(new_n634), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n557), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n450), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n487), .ZN(G1324gat));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n489), .B1(new_n662), .B2(new_n288), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G8gat), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n659), .A2(new_n410), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT42), .B2(new_n666), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n659), .B2(new_n447), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n376), .A2(new_n377), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n484), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n659), .B2(new_n671), .ZN(G1326gat));
  NOR2_X1   g471(.A1(new_n659), .A2(new_n407), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n450), .ZN(new_n676));
  INV_X1    g475(.A(new_n634), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n656), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n595), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT106), .Z(new_n680));
  NAND4_X1  g479(.A1(new_n557), .A2(new_n676), .A3(new_n475), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  INV_X1    g481(.A(new_n594), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n592), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n448), .A2(new_n451), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n450), .A2(new_n402), .A3(new_n410), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n414), .B1(new_n686), .B2(KEYINPUT35), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n452), .A2(KEYINPUT44), .A3(new_n684), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n556), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n450), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n682), .B1(new_n696), .B2(new_n475), .ZN(G1328gat));
  NAND4_X1  g496(.A1(new_n557), .A2(new_n461), .A3(new_n288), .A4(new_n680), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n695), .B2(new_n410), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NOR2_X1   g500(.A1(new_n447), .A2(new_n458), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n692), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n557), .A2(new_n670), .A3(new_n680), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n704), .A2(new_n458), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n705));
  OR2_X1    g504(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n703), .B2(new_n705), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(G1330gat));
  NOR2_X1   g508(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT109), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n690), .A2(new_n401), .A3(new_n691), .A4(new_n694), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n407), .A2(G50gat), .ZN(new_n714));
  AND4_X1   g513(.A1(new_n452), .A2(new_n556), .A3(new_n680), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n715), .B1(new_n712), .B2(G50gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n718), .ZN(new_n721));
  INV_X1    g520(.A(new_n711), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n719), .A2(new_n723), .ZN(G1331gat));
  NOR4_X1   g523(.A1(new_n677), .A2(new_n684), .A3(new_n556), .A4(new_n656), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n452), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n676), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n288), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT49), .B(G64gat), .Z(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(G1333gat));
  INV_X1    g531(.A(new_n447), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n670), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(G71gat), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n734), .A2(G71gat), .B1(new_n726), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n726), .A2(new_n401), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT110), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n556), .A2(new_n634), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n655), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n692), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n450), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n684), .B(new_n742), .C1(new_n685), .C2(new_n687), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT113), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  INV_X1    g551(.A(new_n688), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n742), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n452), .A2(KEYINPUT51), .A3(new_n684), .A4(new_n742), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n750), .A2(new_n752), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n676), .A2(new_n569), .A3(new_n655), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n746), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  NAND4_X1  g559(.A1(new_n690), .A2(new_n288), .A3(new_n691), .A4(new_n744), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(new_n761), .B2(G92gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n288), .A2(new_n570), .A3(new_n655), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT114), .Z(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n747), .A2(KEYINPUT115), .A3(new_n748), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n755), .A2(new_n756), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n755), .A2(new_n756), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n764), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(new_n772), .B1(G92gat), .B2(new_n761), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n765), .B1(new_n773), .B2(new_n774), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n745), .B2(new_n447), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n735), .A2(G99gat), .A3(new_n656), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n758), .B2(new_n777), .ZN(G1338gat));
  NAND4_X1  g577(.A1(new_n690), .A2(new_n401), .A3(new_n691), .A4(new_n744), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n779), .B2(G106gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n407), .A2(G106gat), .A3(new_n656), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n758), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n771), .A2(new_n781), .B1(G106gat), .B2(new_n779), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n657), .A2(new_n556), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n644), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n646), .B1(new_n640), .B2(new_n641), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n651), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n654), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n792), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n453), .B1(new_n530), .B2(new_n524), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n509), .A2(new_n455), .A3(new_n510), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n546), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n554), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n684), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n554), .A2(new_n655), .A3(new_n800), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n556), .B2(new_n797), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(new_n684), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n787), .B1(new_n805), .B2(new_n677), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n401), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n450), .A2(new_n288), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n670), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(new_n293), .A3(new_n693), .ZN(new_n810));
  NOR4_X1   g609(.A1(new_n806), .A2(new_n450), .A3(new_n288), .A4(new_n409), .ZN(new_n811));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n556), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n810), .A2(new_n812), .ZN(G1340gat));
  OAI21_X1  g612(.A(G120gat), .B1(new_n809), .B2(new_n656), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n301), .A3(new_n655), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1341gat));
  OAI21_X1  g615(.A(G127gat), .B1(new_n809), .B2(new_n677), .ZN(new_n817));
  INV_X1    g616(.A(G127gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n818), .A3(new_n634), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n811), .A2(new_n821), .A3(new_n684), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n809), .B2(new_n595), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(G1343gat));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT55), .B1(new_n796), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n789), .A2(KEYINPUT116), .A3(new_n792), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n794), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n555), .A2(new_n554), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n549), .B1(new_n533), .B2(new_n540), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(KEYINPUT94), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n803), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n684), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g635(.A1(new_n594), .A2(new_n593), .A3(new_n797), .A4(new_n801), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n677), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n658), .A2(new_n693), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n841), .B2(new_n407), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n793), .A2(new_n654), .ZN(new_n844));
  INV_X1    g643(.A(new_n796), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(KEYINPUT55), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n541), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(new_n547), .B1(new_n832), .B2(KEYINPUT94), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n553), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n595), .B1(new_n849), .B2(new_n803), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n634), .B1(new_n850), .B2(new_n802), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n843), .B(new_n401), .C1(new_n851), .C2(new_n787), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n808), .A2(new_n447), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n842), .A2(new_n556), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G141gat), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n806), .A2(new_n450), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n733), .A2(new_n407), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n410), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n693), .A2(G141gat), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n855), .B(new_n856), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n859), .A2(new_n288), .A3(new_n864), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(new_n856), .ZN(G1344gat));
  INV_X1    g669(.A(G148gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT59), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n842), .A2(new_n852), .A3(new_n853), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n656), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n401), .A2(new_n843), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n840), .B2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n838), .A2(new_n878), .A3(new_n839), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n401), .B1(new_n851), .B2(new_n787), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n877), .A2(new_n879), .B1(KEYINPUT57), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n808), .A2(new_n447), .A3(new_n655), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n875), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n790), .A3(new_n791), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n642), .A2(new_n791), .A3(new_n643), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n652), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n827), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n795), .A3(new_n829), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n844), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n848), .B2(new_n553), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n595), .B1(new_n891), .B2(new_n803), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n634), .B1(new_n892), .B2(new_n802), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n893), .B2(new_n787), .ZN(new_n894));
  INV_X1    g693(.A(new_n876), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n879), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n806), .B2(new_n407), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n875), .A3(new_n897), .A4(new_n882), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G148gat), .ZN(new_n899));
  OAI211_X1 g698(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n883), .C2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n897), .A3(new_n882), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(G148gat), .A3(new_n898), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT121), .B1(new_n904), .B2(KEYINPUT59), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n874), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n863), .A2(G148gat), .A3(new_n656), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(G155gat), .B1(new_n873), .B2(new_n677), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n677), .A2(G155gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n863), .B2(new_n910), .ZN(G1346gat));
  NAND2_X1  g710(.A1(new_n684), .A2(new_n311), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n873), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n863), .A2(new_n595), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n311), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g716(.A(KEYINPUT122), .B(new_n913), .C1(new_n914), .C2(new_n311), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  NAND2_X1  g718(.A1(new_n450), .A2(new_n288), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n735), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n807), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n807), .A2(KEYINPUT123), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n248), .A3(new_n693), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n806), .A2(new_n676), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n288), .A3(new_n402), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n556), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n927), .A2(new_n931), .ZN(G1348gat));
  OAI21_X1  g731(.A(G176gat), .B1(new_n926), .B2(new_n656), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n249), .A3(new_n655), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n926), .B2(new_n677), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n235), .A3(new_n634), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n930), .A2(new_n234), .A3(new_n684), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n684), .A3(new_n925), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  AND4_X1   g741(.A1(KEYINPUT124), .A2(new_n941), .A3(new_n942), .A4(G190gat), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n226), .B1(new_n944), .B2(KEYINPUT61), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n941), .A2(new_n945), .B1(KEYINPUT124), .B2(new_n942), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n943), .B2(new_n946), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n733), .A2(new_n920), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n881), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(G197gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n949), .A2(new_n950), .A3(new_n693), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n733), .A2(new_n410), .A3(new_n407), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n928), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n556), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(new_n953), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(G204gat), .A3(new_n656), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n949), .B2(new_n656), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n953), .A2(new_n261), .A3(new_n634), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n881), .A2(new_n634), .A3(new_n948), .ZN(new_n963));
  AND4_X1   g762(.A1(new_n962), .A2(new_n963), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n261), .B1(KEYINPUT125), .B2(new_n965), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n963), .A2(new_n966), .B1(new_n962), .B2(KEYINPUT63), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n961), .B1(new_n964), .B2(new_n967), .ZN(G1354gat));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n595), .B1(new_n949), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n969), .B2(new_n949), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G218gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n262), .A3(new_n684), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


