//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT80), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n190), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT79), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n188), .B(KEYINPUT3), .C1(new_n190), .C2(new_n191), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n189), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(new_n192), .B2(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(new_n203), .A3(new_n196), .A4(new_n197), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT4), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT81), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n200), .B(G101), .C1(KEYINPUT81), .C2(new_n205), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n207), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n195), .B2(new_n198), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n204), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(new_n211), .ZN(new_n222));
  OAI211_X1 g036(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n210), .C2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G128), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT64), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n214), .A2(new_n227), .A3(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n232), .B2(new_n214), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n204), .A2(new_n220), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n219), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n243), .A3(new_n246), .A4(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n237), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n219), .A2(new_n230), .A3(new_n250), .A4(new_n236), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G110), .B(G140), .ZN(new_n253));
  INV_X1    g067(.A(G227), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G953), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n253), .B(new_n255), .Z(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n187), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  AOI211_X1 g072(.A(KEYINPUT85), .B(new_n256), .C1(new_n249), .C2(new_n251), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n234), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n229), .B1(new_n204), .B2(new_n220), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT82), .B(new_n248), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT12), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n234), .B1(new_n221), .B2(new_n229), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n265), .A2(KEYINPUT82), .A3(new_n266), .A4(new_n248), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n251), .A2(new_n256), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT72), .B(G902), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT84), .B(G469), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n264), .A2(new_n267), .A3(new_n251), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT83), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n264), .A2(new_n267), .A3(new_n251), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n257), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n249), .A2(new_n256), .A3(new_n251), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G469), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n231), .A2(G119), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G119), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G128), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G110), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT76), .Z(new_n297));
  AND2_X1   g111(.A1(new_n289), .A2(new_n293), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT24), .B(G110), .Z(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G125), .B(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n208), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n301), .B2(KEYINPUT16), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(G146), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n299), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n309), .A2(new_n310), .B1(new_n295), .B2(G110), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n305), .A2(G146), .ZN(new_n312));
  OAI221_X1 g126(.A(new_n311), .B1(new_n310), .B2(new_n309), .C1(new_n306), .C2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT75), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G221), .A3(G234), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(G137), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n308), .A2(new_n314), .A3(new_n320), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n274), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  INV_X1    g139(.A(G217), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n274), .B2(G234), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n322), .A2(new_n328), .A3(new_n274), .A4(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n322), .A2(new_n323), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n327), .A2(G902), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT78), .Z(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT9), .B(G234), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G221), .B1(new_n337), .B2(G902), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n288), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n316), .A2(G952), .ZN(new_n341));
  NAND2_X1  g155(.A1(G234), .A2(G237), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n273), .A2(G953), .A3(new_n342), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT21), .B(G898), .Z(new_n345));
  OAI21_X1  g159(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n346), .B(KEYINPUT94), .Z(new_n347));
  OAI21_X1  g161(.A(G214), .B1(G237), .B2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n350));
  INV_X1    g164(.A(G116), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(G119), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(G119), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n292), .A2(KEYINPUT65), .A3(G116), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G113), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT2), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G113), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n359), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(new_n353), .A3(new_n352), .A4(new_n354), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n207), .A2(new_n364), .A3(new_n218), .ZN(new_n365));
  INV_X1    g179(.A(new_n363), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n355), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n351), .A2(G119), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n356), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n221), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(G110), .B(G122), .Z(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n376), .A3(new_n372), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n222), .A2(KEYINPUT1), .A3(new_n231), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G128), .A3(new_n223), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n222), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n303), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n216), .A2(G125), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n386), .A2(KEYINPUT87), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(KEYINPUT87), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G224), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n389), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n373), .A2(new_n393), .A3(new_n374), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n378), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT7), .ZN(new_n396));
  OR3_X1    g210(.A1(new_n389), .A2(new_n396), .A3(new_n391), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n385), .A2(new_n386), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n396), .B2(new_n391), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n204), .A2(new_n220), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n371), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n374), .B(KEYINPUT8), .Z(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n355), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n366), .B1(new_n404), .B2(new_n370), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n401), .B(new_n402), .C1(new_n400), .C2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n397), .A2(new_n399), .A3(new_n406), .A4(new_n377), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n395), .A2(new_n285), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n409), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n395), .A2(new_n285), .A3(new_n413), .A4(new_n407), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n349), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G475), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(G104), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT19), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT90), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n301), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(G125), .A2(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(G125), .A2(G140), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT90), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n421), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT19), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT91), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n426), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT90), .B1(new_n424), .B2(new_n425), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT19), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n208), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G237), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n316), .A3(G214), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n210), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n436), .A2(new_n316), .A3(G143), .A4(G214), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n246), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n246), .A3(new_n439), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n306), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G146), .B1(new_n430), .B2(new_n431), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n302), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT18), .A2(G131), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n438), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(KEYINPUT89), .A3(KEYINPUT18), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT89), .B1(new_n440), .B2(KEYINPUT18), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n446), .B(new_n449), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n420), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n305), .B(new_n208), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n441), .A2(new_n456), .A3(new_n442), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n455), .B(new_n457), .C1(new_n456), .C2(new_n441), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n458), .A2(new_n453), .A3(new_n420), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n417), .B(new_n285), .C1(new_n454), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT20), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n453), .A3(new_n420), .ZN(new_n462));
  INV_X1    g276(.A(new_n452), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n448), .B1(new_n463), .B2(new_n450), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n464), .A2(new_n446), .B1(new_n435), .B2(new_n443), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n465), .B2(new_n420), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(KEYINPUT92), .C1(G475), .C2(G902), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n468), .A3(new_n417), .A4(new_n285), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n461), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n420), .B1(new_n458), .B2(new_n453), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n285), .B1(new_n459), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G475), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(KEYINPUT92), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G116), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n351), .A2(G122), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n189), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(KEYINPUT14), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G128), .B(G143), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n239), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n481), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n189), .A2(KEYINPUT14), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n484), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(KEYINPUT13), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n210), .A2(G128), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n490), .B(G134), .C1(KEYINPUT13), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n239), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n487), .A2(G107), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n492), .B(new_n493), .C1(new_n494), .C2(new_n482), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n337), .A2(new_n326), .A3(G953), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n274), .ZN(new_n502));
  INV_X1    g316(.A(G478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n502), .B(new_n504), .Z(new_n505));
  NAND2_X1  g319(.A1(new_n476), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n416), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n242), .A2(G134), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n239), .A2(G137), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n247), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n226), .B2(new_n228), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n216), .B1(new_n247), .B2(new_n245), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT30), .ZN(new_n514));
  INV_X1    g328(.A(new_n512), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n248), .A2(new_n516), .A3(new_n217), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n248), .B2(new_n217), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n514), .B1(new_n519), .B2(KEYINPUT30), .ZN(new_n520));
  INV_X1    g334(.A(new_n364), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT67), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n248), .A2(new_n217), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT66), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n513), .A2(new_n516), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n524), .B1(new_n528), .B2(new_n515), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n523), .B(new_n364), .C1(new_n529), .C2(new_n514), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n361), .A2(new_n363), .A3(KEYINPUT68), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT68), .B1(new_n361), .B2(new_n363), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n436), .A2(new_n316), .A3(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n203), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n538), .B(new_n539), .Z(new_n540));
  NAND4_X1  g354(.A1(new_n531), .A2(new_n532), .A3(new_n536), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT69), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n525), .B(new_n542), .C1(new_n384), .C2(new_n511), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT69), .B1(new_n512), .B2(new_n513), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n535), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n364), .B1(new_n512), .B2(new_n513), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n536), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n540), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n522), .A2(new_n530), .A3(new_n536), .A4(new_n540), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n541), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT32), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G472), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n522), .A2(new_n530), .A3(new_n536), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n555), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n550), .A2(new_n565), .A3(new_n553), .A4(new_n540), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n545), .A2(new_n547), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT70), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n568), .A2(new_n553), .A3(new_n569), .A4(new_n540), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT71), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n564), .A2(new_n566), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n519), .B1(new_n533), .B2(new_n534), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n536), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT28), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n550), .A2(KEYINPUT29), .A3(new_n540), .A4(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(new_n274), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n562), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n561), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n559), .A2(KEYINPUT32), .A3(new_n560), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT73), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT73), .ZN(new_n584));
  NOR4_X1   g398(.A1(new_n583), .A2(new_n561), .A3(new_n579), .A4(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n340), .B(new_n507), .C1(new_n582), .C2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND2_X1  g401(.A1(new_n408), .A2(new_n410), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n395), .A2(new_n285), .A3(new_n411), .A4(new_n407), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n348), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n347), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n461), .A2(new_n467), .A3(new_n469), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n473), .C1(new_n469), .C2(new_n474), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n501), .A2(KEYINPUT33), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n499), .B2(new_n500), .ZN(new_n597));
  OAI211_X1 g411(.A(G478), .B(new_n274), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n502), .A2(new_n503), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT95), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n562), .B1(new_n559), .B2(new_n274), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n559), .A2(new_n560), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n603), .A2(new_n339), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NOR2_X1   g424(.A1(new_n339), .A2(new_n607), .ZN(new_n611));
  INV_X1    g425(.A(new_n505), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n461), .A2(new_n469), .B1(G475), .B2(new_n472), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n592), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NOR2_X1   g433(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n315), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n333), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n330), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n258), .A2(new_n259), .A3(new_n270), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n624), .A2(new_n273), .A3(new_n275), .ZN(new_n625));
  INV_X1    g439(.A(G469), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n284), .B2(new_n285), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n338), .B(new_n623), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n507), .A3(new_n606), .A4(new_n605), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  OAI21_X1  g446(.A(new_n343), .B1(new_n344), .B2(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n614), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n591), .B(new_n635), .C1(new_n582), .C2(new_n585), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  INV_X1    g451(.A(KEYINPUT32), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n606), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n563), .A2(new_n540), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n640), .B(new_n285), .C1(new_n540), .C2(new_n575), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G472), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n639), .A2(new_n581), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT97), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n612), .A2(new_n594), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n412), .A2(new_n414), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT96), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT38), .ZN(new_n649));
  INV_X1    g463(.A(new_n348), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n650), .A3(new_n623), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n288), .A2(new_n338), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n633), .B(KEYINPUT39), .Z(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT98), .Z(new_n655));
  AND2_X1   g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n646), .B(new_n651), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G143), .ZN(G45));
  OAI211_X1 g473(.A(new_n600), .B(new_n633), .C1(new_n470), .C2(new_n475), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n590), .A2(new_n660), .A3(KEYINPUT99), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n628), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT99), .B1(new_n590), .B2(new_n660), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n662), .B(new_n663), .C1(new_n582), .C2(new_n585), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n573), .A2(new_n578), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n639), .A2(new_n581), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n584), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n580), .A2(KEYINPUT73), .A3(new_n581), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(KEYINPUT100), .A3(new_n662), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT101), .B(G146), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G48));
  OAI21_X1  g491(.A(G469), .B1(new_n624), .B2(new_n273), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n277), .A2(new_n678), .A3(new_n338), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n671), .A2(new_n672), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n335), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n603), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT41), .B(G113), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NOR3_X1   g500(.A1(new_n683), .A2(new_n592), .A3(new_n615), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n351), .ZN(G18));
  INV_X1    g502(.A(new_n506), .ZN(new_n689));
  INV_X1    g503(.A(new_n623), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n679), .A2(new_n590), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n682), .A2(new_n689), .A3(new_n347), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  INV_X1    g507(.A(new_n645), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n681), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n335), .B(KEYINPUT105), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n605), .A2(KEYINPUT104), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT104), .B(new_n562), .C1(new_n559), .C2(new_n274), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n560), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n557), .B(new_n532), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n550), .A2(new_n576), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n555), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT103), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n707), .B(new_n701), .C1(new_n702), .C2(new_n704), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n698), .A2(new_n700), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n696), .B1(new_n697), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  OAI22_X1  g526(.A1(new_n604), .A2(new_n712), .B1(new_n705), .B2(KEYINPUT103), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n708), .A3(new_n699), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n335), .B(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(KEYINPUT106), .A3(new_n715), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n592), .B(new_n695), .C1(new_n711), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n477), .ZN(G24));
  NOR2_X1   g532(.A1(new_n713), .A2(new_n699), .ZN(new_n719));
  INV_X1    g533(.A(new_n660), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n691), .A3(new_n720), .A4(new_n709), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  XOR2_X1   g536(.A(new_n581), .B(KEYINPUT107), .Z(new_n723));
  AOI21_X1  g537(.A(new_n697), .B1(new_n580), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n647), .A2(new_n660), .A3(new_n650), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT42), .B1(new_n726), .B2(new_n652), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n339), .B1(new_n671), .B2(new_n672), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n647), .A2(new_n650), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  INV_X1    g547(.A(new_n634), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n728), .A2(new_n734), .A3(new_n729), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  XNOR2_X1  g550(.A(new_n284), .B(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(G469), .C1(new_n737), .C2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n277), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n338), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n653), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n476), .A2(new_n600), .ZN(new_n746));
  NAND2_X1  g560(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n476), .A2(new_n600), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n607), .A3(new_n623), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n745), .B1(KEYINPUT44), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n729), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n242), .ZN(G39));
  OR2_X1    g572(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n744), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n744), .A2(new_n759), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n682), .A2(new_n335), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n725), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n770));
  INV_X1    g584(.A(new_n679), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n729), .ZN(new_n772));
  INV_X1    g586(.A(new_n343), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n751), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT118), .Z(new_n776));
  INV_X1    g590(.A(new_n724), .ZN(new_n777));
  OR4_X1    g591(.A1(new_n770), .A2(new_n776), .A3(KEYINPUT48), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n770), .A2(KEYINPUT48), .ZN(new_n779));
  OAI22_X1  g593(.A1(new_n776), .A2(new_n777), .B1(new_n770), .B2(KEYINPUT48), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n772), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n644), .A2(new_n773), .A3(new_n335), .A4(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n781), .B(new_n341), .C1(new_n601), .C2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n594), .A3(new_n600), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n776), .A2(new_n690), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(new_n714), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n774), .B1(new_n711), .B2(new_n716), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n650), .A3(new_n649), .A4(new_n771), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT50), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n277), .A2(new_n678), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n338), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n729), .B(new_n788), .C1(new_n763), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n789), .A2(new_n791), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n787), .A2(new_n792), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT51), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n784), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n788), .A2(new_n591), .A3(new_n771), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n590), .B1(new_n671), .B2(new_n672), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n713), .A2(new_n660), .A3(new_n699), .A4(new_n708), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n806), .A2(new_n635), .B1(new_n807), .B2(new_n691), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n633), .B(KEYINPUT114), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n652), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n645), .A2(new_n590), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n690), .A3(new_n643), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n664), .A2(new_n665), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT100), .B1(new_n673), .B2(new_n662), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n808), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n636), .A2(new_n721), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n666), .B2(new_n674), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .A3(new_n812), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n629), .A2(new_n729), .ZN(new_n822));
  INV_X1    g636(.A(new_n633), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n612), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n613), .B(new_n824), .C1(new_n582), .C2(new_n585), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n714), .A2(new_n720), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n682), .A2(new_n340), .A3(new_n734), .A4(new_n729), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT113), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  INV_X1    g644(.A(new_n824), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n671), .B2(new_n672), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n807), .B1(new_n832), .B2(new_n613), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n830), .B(new_n735), .C1(new_n833), .C2(new_n822), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n594), .A2(new_n505), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n415), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n415), .B2(new_n836), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n837), .A2(new_n838), .B1(new_n416), .B2(new_n601), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n611), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n586), .A2(new_n840), .A3(new_n841), .A4(new_n630), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n586), .A2(new_n840), .A3(new_n630), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT112), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n829), .A2(new_n834), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n692), .B1(new_n603), .B2(new_n683), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n717), .A2(new_n687), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n821), .A2(new_n732), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(new_n819), .B2(new_n812), .ZN(new_n853));
  AND4_X1   g667(.A1(KEYINPUT52), .A2(new_n675), .A3(new_n808), .A4(new_n812), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n845), .B(KEYINPUT115), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n848), .B1(KEYINPUT53), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n804), .A2(new_n805), .A3(new_n851), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(G952), .B2(G953), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n649), .A2(new_n338), .A3(new_n715), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n793), .B(KEYINPUT49), .Z(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n746), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n861), .A2(new_n348), .A3(new_n863), .A4(new_n644), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(G75));
  INV_X1    g679(.A(new_n848), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n855), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n273), .A3(new_n411), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT120), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n378), .A2(new_n394), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(new_n392), .Z(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n875), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n316), .A2(G952), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G51));
  XOR2_X1   g693(.A(new_n739), .B(KEYINPUT57), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n856), .A2(new_n857), .A3(new_n852), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT54), .B1(new_n868), .B2(new_n869), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n272), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n856), .A2(new_n857), .A3(new_n274), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(G469), .A3(new_n737), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n878), .B1(new_n884), .B2(new_n886), .ZN(G54));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(KEYINPUT58), .B2(G475), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n466), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n878), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n885), .A2(new_n466), .A3(new_n890), .A4(new_n891), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G60));
  NOR2_X1   g711(.A1(new_n595), .A2(new_n597), .ZN(new_n898));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n881), .B2(new_n882), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n851), .B2(new_n858), .ZN(new_n903));
  INV_X1    g717(.A(new_n898), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n902), .B(new_n895), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(G63));
  NOR2_X1   g720(.A1(new_n856), .A2(new_n857), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT60), .Z(new_n909));
  NAND4_X1  g723(.A1(new_n907), .A2(KEYINPUT122), .A3(new_n621), .A4(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n868), .A2(new_n869), .A3(new_n909), .ZN(new_n911));
  INV_X1    g725(.A(new_n331), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n878), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n868), .A2(new_n621), .A3(new_n869), .A4(new_n909), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n910), .A2(new_n913), .A3(KEYINPUT61), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G66));
  INV_X1    g735(.A(new_n345), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n922), .B2(new_n390), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n844), .A2(new_n842), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n847), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n847), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n873), .B1(G898), .B2(new_n316), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  INV_X1    g745(.A(new_n732), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n766), .B2(new_n767), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n745), .A2(new_n724), .A3(new_n811), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT124), .Z(new_n935));
  INV_X1    g749(.A(new_n757), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n936), .A2(new_n735), .A3(new_n819), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n429), .A2(new_n434), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n520), .B(new_n939), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n601), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n655), .B(new_n729), .C1(new_n943), .C2(new_n836), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n682), .A2(new_n335), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n766), .B2(new_n767), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n658), .A2(KEYINPUT62), .A3(new_n819), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT62), .B1(new_n658), .B2(new_n819), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n947), .B(new_n936), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n942), .B(new_n316), .C1(new_n941), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n940), .B1(KEYINPUT125), .B2(G900), .ZN(new_n952));
  AND2_X1   g766(.A1(G227), .A2(G900), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n952), .B(new_n954), .C1(KEYINPUT125), .C2(G900), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n955), .B(G953), .C1(new_n941), .C2(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n951), .A2(new_n956), .ZN(G72));
  NAND4_X1  g771(.A1(new_n933), .A2(new_n555), .A3(new_n935), .A4(new_n937), .ZN(new_n958));
  OAI22_X1  g772(.A1(new_n950), .A2(new_n640), .B1(new_n958), .B2(new_n563), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n878), .B1(new_n959), .B2(new_n928), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n564), .A2(new_n557), .ZN(new_n961));
  XNOR2_X1  g775(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n562), .A2(new_n285), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n850), .A2(new_n961), .A3(new_n964), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(G57));
endmodule


