

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n722), .ZN(n707) );
  NAND2_X1 U551 ( .A1(G8), .A2(n722), .ZN(n772) );
  AND2_X2 U552 ( .A1(n522), .A2(G2104), .ZN(n888) );
  INV_X1 U553 ( .A(KEYINPUT97), .ZN(n699) );
  NAND2_X1 U554 ( .A1(n517), .A2(n516), .ZN(n807) );
  AND2_X1 U555 ( .A1(n525), .A2(n514), .ZN(G164) );
  AND2_X1 U556 ( .A1(n524), .A2(n523), .ZN(n514) );
  AND2_X1 U557 ( .A1(n982), .A2(n817), .ZN(n515) );
  OR2_X1 U558 ( .A1(n772), .A2(n771), .ZN(n516) );
  AND2_X1 U559 ( .A1(n769), .A2(n768), .ZN(n517) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n685) );
  NOR2_X1 U561 ( .A1(n805), .A2(n515), .ZN(n806) );
  XNOR2_X1 U562 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n540) );
  NOR2_X2 U563 ( .A1(n613), .A2(n542), .ZN(n641) );
  NOR2_X1 U564 ( .A1(G651), .A2(n613), .ZN(n642) );
  XNOR2_X1 U565 ( .A(n541), .B(n540), .ZN(n550) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT87), .ZN(n525) );
  XNOR2_X1 U567 ( .A(KEYINPUT7), .B(n551), .ZN(G168) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n522), .ZN(n883) );
  NAND2_X1 U569 ( .A1(G126), .A2(n883), .ZN(n519) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U571 ( .A1(G114), .A2(n884), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U574 ( .A(KEYINPUT17), .B(n521), .Z(n531) );
  NAND2_X1 U575 ( .A1(G138), .A2(n531), .ZN(n524) );
  INV_X1 U576 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U577 ( .A1(G102), .A2(n888), .ZN(n523) );
  INV_X1 U578 ( .A(KEYINPUT65), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n888), .A2(G101), .ZN(n526) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n526), .Z(n528) );
  NAND2_X1 U581 ( .A1(n883), .A2(G125), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U583 ( .A(n530), .B(n529), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G113), .A2(n884), .ZN(n533) );
  BUF_X1 U585 ( .A(n531), .Z(n887) );
  NAND2_X1 U586 ( .A1(G137), .A2(n887), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U588 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U590 ( .A1(n637), .A2(G89), .ZN(n536) );
  XOR2_X1 U591 ( .A(KEYINPUT4), .B(n536), .Z(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n613) );
  INV_X1 U593 ( .A(G651), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n641), .A2(G76), .ZN(n537) );
  XOR2_X1 U595 ( .A(KEYINPUT76), .B(n537), .Z(n538) );
  NOR2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n642), .A2(G51), .ZN(n546) );
  NOR2_X1 U598 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n543), .Z(n544) );
  XNOR2_X1 U600 ( .A(KEYINPUT66), .B(n544), .ZN(n638) );
  NAND2_X1 U601 ( .A1(G63), .A2(n638), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n548) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n547) );
  XNOR2_X1 U604 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n551) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U607 ( .A1(G123), .A2(n883), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT18), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G111), .A2(n884), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G135), .A2(n887), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G99), .A2(n888), .ZN(n555) );
  XNOR2_X1 U613 ( .A(KEYINPUT79), .B(n555), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n930) );
  XNOR2_X1 U616 ( .A(G2096), .B(n930), .ZN(n560) );
  OR2_X1 U617 ( .A1(G2100), .A2(n560), .ZN(G156) );
  INV_X1 U618 ( .A(G132), .ZN(G219) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  NAND2_X1 U621 ( .A1(G90), .A2(n637), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G77), .A2(n641), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT9), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G52), .A2(n642), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G64), .A2(n638), .ZN(n566) );
  XNOR2_X1 U628 ( .A(KEYINPUT69), .B(n566), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(G171) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT72), .ZN(n570) );
  XNOR2_X1 U633 ( .A(KEYINPUT10), .B(n570), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n833) );
  NAND2_X1 U635 ( .A1(n833), .A2(G567), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT11), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT73), .B(n572), .ZN(G234) );
  INV_X1 U638 ( .A(G860), .ZN(n840) );
  XNOR2_X1 U639 ( .A(KEYINPUT74), .B(n840), .ZN(n602) );
  NAND2_X1 U640 ( .A1(n638), .A2(G56), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n573), .Z(n579) );
  NAND2_X1 U642 ( .A1(n637), .A2(G81), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G68), .A2(n641), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n642), .A2(G43), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n990) );
  OR2_X1 U650 ( .A1(n602), .A2(n990), .ZN(G153) );
  INV_X1 U651 ( .A(G171), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G92), .A2(n637), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G66), .A2(n638), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U655 ( .A1(G79), .A2(n641), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G54), .A2(n642), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n588), .Z(n977) );
  NOR2_X1 U660 ( .A1(n977), .A2(G868), .ZN(n589) );
  XNOR2_X1 U661 ( .A(n589), .B(KEYINPUT75), .ZN(n591) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n637), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G78), .A2(n641), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U667 ( .A(KEYINPUT70), .B(n594), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G53), .A2(n642), .ZN(n595) );
  XNOR2_X1 U669 ( .A(KEYINPUT71), .B(n595), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G65), .A2(n638), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(G299) );
  INV_X1 U673 ( .A(G868), .ZN(n657) );
  NOR2_X1 U674 ( .A1(G286), .A2(n657), .ZN(n601) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n603), .A2(n977), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n990), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G868), .A2(n977), .ZN(n605) );
  NOR2_X1 U682 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G74), .A2(G651), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT82), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G49), .A2(n642), .ZN(n609) );
  XOR2_X1 U687 ( .A(KEYINPUT81), .B(n609), .Z(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n638), .A2(n612), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n613), .A2(G87), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G288) );
  NAND2_X1 U692 ( .A1(G88), .A2(n637), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G75), .A2(n641), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n642), .A2(G50), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G62), .A2(n638), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(G166) );
  NAND2_X1 U699 ( .A1(n642), .A2(G47), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT68), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G85), .A2(n637), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G72), .A2(n641), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G60), .A2(n638), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT67), .B(n625), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G290) );
  NAND2_X1 U708 ( .A1(G86), .A2(n637), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G61), .A2(n638), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n641), .A2(G73), .ZN(n632) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n642), .A2(G48), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G93), .A2(n637), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G67), .A2(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n646) );
  NAND2_X1 U719 ( .A1(G80), .A2(n641), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G55), .A2(n642), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U723 ( .A(KEYINPUT80), .B(n647), .Z(n843) );
  XNOR2_X1 U724 ( .A(G166), .B(KEYINPUT19), .ZN(n649) );
  INV_X1 U725 ( .A(G299), .ZN(n681) );
  XNOR2_X1 U726 ( .A(G290), .B(n681), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U728 ( .A(n650), .B(G305), .Z(n651) );
  XNOR2_X1 U729 ( .A(G288), .B(n651), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n843), .B(n652), .ZN(n911) );
  NAND2_X1 U731 ( .A1(G559), .A2(n977), .ZN(n653) );
  XOR2_X1 U732 ( .A(n990), .B(n653), .Z(n841) );
  XNOR2_X1 U733 ( .A(n911), .B(n841), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n654), .B(KEYINPUT83), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n655), .A2(G868), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT84), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n843), .A2(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G2072), .ZN(n664) );
  XOR2_X1 U744 ( .A(KEYINPUT85), .B(n664), .Z(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U746 ( .A1(G120), .A2(G69), .ZN(n665) );
  NOR2_X1 U747 ( .A1(G237), .A2(n665), .ZN(n666) );
  XNOR2_X1 U748 ( .A(KEYINPUT86), .B(n666), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n667), .A2(G108), .ZN(n844) );
  NAND2_X1 U750 ( .A1(G567), .A2(n844), .ZN(n672) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U753 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G96), .A2(n670), .ZN(n845) );
  NAND2_X1 U755 ( .A1(G2106), .A2(n845), .ZN(n671) );
  NAND2_X1 U756 ( .A1(n672), .A2(n671), .ZN(n846) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U758 ( .A1(n846), .A2(n673), .ZN(n839) );
  NAND2_X1 U759 ( .A1(n839), .A2(G36), .ZN(G176) );
  XOR2_X1 U760 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n789) );
  INV_X1 U762 ( .A(n789), .ZN(n674) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n790) );
  NAND2_X2 U764 ( .A1(n674), .A2(n790), .ZN(n722) );
  NAND2_X1 U765 ( .A1(n707), .A2(G2072), .ZN(n675) );
  XNOR2_X1 U766 ( .A(n675), .B(KEYINPUT27), .ZN(n677) );
  INV_X1 U767 ( .A(G1956), .ZN(n1005) );
  NOR2_X1 U768 ( .A1(n1005), .A2(n707), .ZN(n676) );
  NOR2_X1 U769 ( .A1(n677), .A2(n676), .ZN(n680) );
  NOR2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n679) );
  INV_X1 U771 ( .A(KEYINPUT28), .ZN(n678) );
  XNOR2_X1 U772 ( .A(n679), .B(n678), .ZN(n691) );
  INV_X1 U773 ( .A(n691), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n681), .A2(n680), .ZN(n682) );
  OR2_X1 U775 ( .A1(n683), .A2(n682), .ZN(n704) );
  INV_X1 U776 ( .A(G1996), .ZN(n684) );
  NOR2_X1 U777 ( .A1(n722), .A2(n684), .ZN(n686) );
  XNOR2_X1 U778 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n722), .A2(G1341), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U781 ( .A1(n990), .A2(n689), .ZN(n696) );
  OR2_X1 U782 ( .A1(n977), .A2(n696), .ZN(n690) );
  AND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n702) );
  NAND2_X1 U784 ( .A1(G1348), .A2(n722), .ZN(n692) );
  XOR2_X1 U785 ( .A(KEYINPUT95), .B(n692), .Z(n695) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n707), .ZN(n693) );
  XNOR2_X1 U787 ( .A(KEYINPUT96), .B(n693), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n696), .A2(n977), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U794 ( .A(KEYINPUT29), .B(n705), .Z(n742) );
  NAND2_X1 U795 ( .A1(G1961), .A2(n722), .ZN(n709) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT94), .Z(n706) );
  XNOR2_X1 U797 ( .A(KEYINPUT25), .B(n706), .ZN(n959) );
  NAND2_X1 U798 ( .A1(n707), .A2(n959), .ZN(n708) );
  NAND2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n720) );
  OR2_X1 U800 ( .A1(G301), .A2(n720), .ZN(n740) );
  INV_X1 U801 ( .A(KEYINPUT99), .ZN(n711) );
  NOR2_X1 U802 ( .A1(G1971), .A2(n772), .ZN(n710) );
  XNOR2_X1 U803 ( .A(n711), .B(n710), .ZN(n713) );
  NOR2_X1 U804 ( .A1(G2090), .A2(n722), .ZN(n712) );
  NOR2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U806 ( .A(KEYINPUT100), .B(n714), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n715), .A2(G303), .ZN(n729) );
  INV_X1 U808 ( .A(n729), .ZN(n716) );
  OR2_X1 U809 ( .A1(n716), .A2(G286), .ZN(n717) );
  AND2_X1 U810 ( .A1(n717), .A2(G8), .ZN(n719) );
  AND2_X1 U811 ( .A1(n740), .A2(n719), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n742), .A2(n718), .ZN(n733) );
  INV_X1 U813 ( .A(n719), .ZN(n731) );
  NAND2_X1 U814 ( .A1(G301), .A2(n720), .ZN(n721) );
  XOR2_X1 U815 ( .A(KEYINPUT98), .B(n721), .Z(n727) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n772), .ZN(n737) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n722), .ZN(n736) );
  NOR2_X1 U818 ( .A1(n737), .A2(n736), .ZN(n723) );
  NAND2_X1 U819 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n725), .A2(G168), .ZN(n726) );
  NOR2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(n728), .Z(n743) );
  AND2_X1 U824 ( .A1(n743), .A2(n729), .ZN(n730) );
  OR2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n735) );
  XOR2_X1 U827 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n734) );
  XNOR2_X1 U828 ( .A(n735), .B(n734), .ZN(n748) );
  AND2_X1 U829 ( .A1(G8), .A2(n736), .ZN(n738) );
  OR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n744) );
  INV_X1 U831 ( .A(n744), .ZN(n739) );
  AND2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n746) );
  OR2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n765) );
  NOR2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n749) );
  XNOR2_X1 U838 ( .A(n749), .B(KEYINPUT102), .ZN(n758) );
  NOR2_X1 U839 ( .A1(G303), .A2(G1971), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n758), .A2(n750), .ZN(n988) );
  NAND2_X1 U841 ( .A1(n765), .A2(n988), .ZN(n751) );
  XNOR2_X1 U842 ( .A(KEYINPUT103), .B(n751), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n976) );
  INV_X1 U844 ( .A(n772), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n976), .A2(n752), .ZN(n753) );
  NOR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U847 ( .A(n755), .B(KEYINPUT64), .ZN(n756) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n756), .ZN(n757) );
  XNOR2_X1 U849 ( .A(G1981), .B(G305), .ZN(n973) );
  NOR2_X1 U850 ( .A1(n757), .A2(n973), .ZN(n762) );
  INV_X1 U851 ( .A(n758), .ZN(n759) );
  NOR2_X1 U852 ( .A1(n772), .A2(n759), .ZN(n760) );
  NAND2_X1 U853 ( .A1(KEYINPUT33), .A2(n760), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G303), .A2(G2090), .ZN(n763) );
  XNOR2_X1 U856 ( .A(KEYINPUT104), .B(n763), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n764), .A2(G8), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n767), .A2(n772), .ZN(n768) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XOR2_X1 U861 ( .A(n770), .B(KEYINPUT24), .Z(n771) );
  NAND2_X1 U862 ( .A1(G119), .A2(n883), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G107), .A2(n884), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G131), .A2(n887), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G95), .A2(n888), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n895) );
  AND2_X1 U869 ( .A1(n895), .A2(G1991), .ZN(n788) );
  NAND2_X1 U870 ( .A1(G105), .A2(n888), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT38), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G117), .A2(n884), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G141), .A2(n887), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G129), .A2(n883), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT91), .B(n782), .ZN(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n901) );
  AND2_X1 U879 ( .A1(n901), .A2(G1996), .ZN(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n935) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n817) );
  INV_X1 U882 ( .A(n817), .ZN(n791) );
  NOR2_X1 U883 ( .A1(n935), .A2(n791), .ZN(n810) );
  XOR2_X1 U884 ( .A(KEYINPUT92), .B(n810), .Z(n803) );
  XNOR2_X1 U885 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NAND2_X1 U886 ( .A1(G140), .A2(n887), .ZN(n793) );
  NAND2_X1 U887 ( .A1(G104), .A2(n888), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n794), .ZN(n801) );
  XNOR2_X1 U890 ( .A(KEYINPUT35), .B(KEYINPUT90), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n883), .A2(G128), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n884), .A2(G116), .ZN(n795) );
  XOR2_X1 U893 ( .A(KEYINPUT89), .B(n795), .Z(n796) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U895 ( .A(n799), .B(n798), .Z(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U897 ( .A(KEYINPUT36), .B(n802), .ZN(n908) );
  NOR2_X1 U898 ( .A1(n815), .A2(n908), .ZN(n922) );
  NAND2_X1 U899 ( .A1(n817), .A2(n922), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n803), .A2(n813), .ZN(n804) );
  XOR2_X1 U901 ( .A(KEYINPUT93), .B(n804), .Z(n805) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n820) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n901), .ZN(n938) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n895), .ZN(n933) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n933), .A2(n808), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n938), .A2(n811), .ZN(n812) );
  XNOR2_X1 U910 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n815), .A2(n908), .ZN(n924) );
  NAND2_X1 U913 ( .A1(n816), .A2(n924), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n822) );
  XOR2_X1 U916 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n821) );
  XNOR2_X1 U917 ( .A(n822), .B(n821), .ZN(G329) );
  XNOR2_X1 U918 ( .A(G2454), .B(G2451), .ZN(n831) );
  XNOR2_X1 U919 ( .A(G2430), .B(G2446), .ZN(n829) );
  XOR2_X1 U920 ( .A(G2435), .B(G2427), .Z(n824) );
  XNOR2_X1 U921 ( .A(KEYINPUT106), .B(G2438), .ZN(n823) );
  XNOR2_X1 U922 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U923 ( .A(n825), .B(G2443), .Z(n827) );
  XNOR2_X1 U924 ( .A(G1341), .B(G1348), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n832), .A2(G14), .ZN(n916) );
  XNOR2_X1 U929 ( .A(KEYINPUT107), .B(n916), .ZN(G401) );
  NAND2_X1 U930 ( .A1(n833), .A2(G2106), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT108), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n836) );
  INV_X1 U933 ( .A(G661), .ZN(n835) );
  NOR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n837), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U938 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  NAND2_X1 U940 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G145) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G108), .ZN(G238) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U947 ( .A(KEYINPUT111), .B(n846), .ZN(G319) );
  XNOR2_X1 U948 ( .A(G1981), .B(G2474), .ZN(n856) );
  XOR2_X1 U949 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1956), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U952 ( .A(G1961), .B(G1986), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U956 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U959 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U962 ( .A(KEYINPUT43), .B(G2090), .Z(n860) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U966 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U968 ( .A1(G124), .A2(n883), .ZN(n865) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n865), .Z(n866) );
  XNOR2_X1 U970 ( .A(n866), .B(KEYINPUT113), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G112), .A2(n884), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G136), .A2(n887), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G100), .A2(n888), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U977 ( .A(KEYINPUT114), .B(n873), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G139), .A2(n887), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G103), .A2(n888), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n882) );
  XNOR2_X1 U981 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n884), .A2(G115), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n883), .A2(G127), .ZN(n876) );
  XOR2_X1 U984 ( .A(KEYINPUT115), .B(n876), .Z(n877) );
  NAND2_X1 U985 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U986 ( .A(n880), .B(n879), .Z(n881) );
  NOR2_X1 U987 ( .A1(n882), .A2(n881), .ZN(n926) );
  NAND2_X1 U988 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U989 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U990 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G142), .A2(n887), .ZN(n890) );
  NAND2_X1 U992 ( .A1(G106), .A2(n888), .ZN(n889) );
  NAND2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  NOR2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n926), .B(n894), .ZN(n907) );
  XNOR2_X1 U997 ( .A(G164), .B(G160), .ZN(n896) );
  XOR2_X1 U998 ( .A(n896), .B(n895), .Z(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT117), .B(KEYINPUT48), .Z(n898) );
  XNOR2_X1 U1000 ( .A(KEYINPUT46), .B(KEYINPUT119), .ZN(n897) );
  XNOR2_X1 U1001 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1002 ( .A(n900), .B(n899), .Z(n905) );
  XOR2_X1 U1003 ( .A(n901), .B(G162), .Z(n902) );
  XNOR2_X1 U1004 ( .A(n902), .B(n930), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n903), .B(KEYINPUT118), .ZN(n904) );
  XNOR2_X1 U1006 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1010 ( .A(n911), .B(G286), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G171), .B(n977), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(n990), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n915), .ZN(G397) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n916), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n922), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n946) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT122), .B(n925), .ZN(n928) );
  XOR2_X1 U1026 ( .A(G2072), .B(n926), .Z(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT50), .B(n929), .ZN(n944) );
  XNOR2_X1 U1029 ( .A(G160), .B(G2084), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT51), .B(KEYINPUT121), .ZN(n940) );
  XOR2_X1 U1034 ( .A(G2090), .B(KEYINPUT120), .Z(n936) );
  XNOR2_X1 U1035 ( .A(G162), .B(n936), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(n940), .B(n939), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1048 ( .A(G2067), .B(G26), .Z(n953) );
  NAND2_X1 U1049 ( .A1(n953), .A2(G28), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G25), .B(G1991), .Z(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT123), .B(n954), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(G27), .B(n959), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT53), .B(n962), .Z(n965) );
  XOR2_X1 U1057 ( .A(KEYINPUT54), .B(G34), .Z(n963) );
  XNOR2_X1 U1058 ( .A(G2084), .B(n963), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1062 ( .A(KEYINPUT55), .B(n968), .Z(n969) );
  NOR2_X1 U1063 ( .A1(G29), .A2(n969), .ZN(n970) );
  XOR2_X1 U1064 ( .A(KEYINPUT124), .B(n970), .Z(n971) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n971), .ZN(n1024) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XOR2_X1 U1067 ( .A(G168), .B(G1966), .Z(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1069 ( .A(KEYINPUT57), .B(n974), .Z(n994) );
  NAND2_X1 U1070 ( .A1(G303), .A2(G1971), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n986) );
  XNOR2_X1 U1072 ( .A(n977), .B(G1348), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n980), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(G1956), .B(G299), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT126), .B(n989), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n990), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1022) );
  INV_X1 U1086 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1087 ( .A(G1966), .B(G21), .Z(n1004) );
  XNOR2_X1 U1088 ( .A(G1986), .B(G24), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(G23), .B(G1976), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT127), .B(n999), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1017) );
  XOR2_X1 U1096 ( .A(G1961), .B(G5), .Z(n1015) );
  XNOR2_X1 U1097 ( .A(G20), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1007) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT59), .B(G1348), .Z(n1010) );
  XNOR2_X1 U1103 ( .A(G4), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(n1013), .B(KEYINPUT60), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

