//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AND4_X1   g018(.A1(new_n200), .A2(new_n202), .A3(new_n204), .A4(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n202), .A2(KEYINPUT77), .A3(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G128), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(new_n204), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n213));
  XNOR2_X1  g027(.A(G104), .B(G107), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G107), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n218), .A2(new_n221), .A3(new_n215), .A4(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n217), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n220), .A2(G104), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT76), .B(G101), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n212), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n206), .A2(G128), .B1(new_n202), .B2(new_n204), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n205), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n199), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT10), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n212), .B2(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n211), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G143), .B(G146), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G128), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT64), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n211), .A2(new_n244), .A3(new_n245), .A4(new_n239), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n240), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G101), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n254), .A2(new_n255), .B1(G131), .B2(new_n193), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n216), .A2(new_n226), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n200), .B1(G143), .B2(new_n201), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n211), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n241), .A2(new_n200), .A3(G128), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n237), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n262), .A3(new_n223), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n238), .A2(new_n253), .A3(new_n256), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n227), .A2(new_n230), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n227), .B2(new_n212), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n266), .A2(KEYINPUT78), .A3(new_n233), .A4(new_n199), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n236), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G227), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT75), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n238), .A2(new_n253), .A3(new_n263), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n238), .A2(new_n253), .A3(KEYINPUT80), .A4(new_n263), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n199), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT79), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n264), .A2(new_n281), .A3(new_n273), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n264), .B2(new_n273), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n275), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G469), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT81), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n264), .A2(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT79), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n264), .A2(new_n281), .A3(new_n273), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n292), .A2(new_n280), .B1(new_n274), .B2(new_n268), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n288), .B(G469), .C1(new_n293), .C2(G902), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT82), .B(G469), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n236), .A2(new_n267), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n264), .A2(new_n298), .A3(new_n273), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n264), .B2(new_n273), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n273), .B1(new_n280), .B2(new_n264), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n295), .B(new_n296), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  OAI21_X1  g119(.A(G221), .B1(new_n305), .B2(G902), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT74), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n243), .A2(new_n246), .ZN(new_n311));
  INV_X1    g125(.A(new_n240), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT84), .B1(new_n247), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n230), .A2(new_n316), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT85), .B(G224), .Z(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G953), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n321), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n315), .A2(new_n317), .A3(new_n323), .A4(new_n318), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT68), .A2(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT68), .A2(G116), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(G119), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G116), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT2), .B(G113), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n332), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n328), .A3(new_n330), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n252), .A3(new_n250), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n330), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n330), .A2(KEYINPUT5), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(G113), .A3(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n257), .A2(new_n340), .A3(new_n335), .A4(new_n223), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G122), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n345), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n341), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT6), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n325), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(G113), .B1(new_n330), .B2(KEYINPUT5), .ZN(new_n351));
  INV_X1    g165(.A(new_n330), .ZN(new_n352));
  INV_X1    g166(.A(new_n327), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT68), .A2(G116), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n355), .B2(G119), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n351), .B1(new_n356), .B2(KEYINPUT5), .ZN(new_n357));
  INV_X1    g171(.A(new_n335), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n227), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n341), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n344), .B(KEYINPUT8), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n319), .A2(new_n321), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n247), .A2(new_n316), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n363), .A2(new_n314), .B1(new_n316), .B2(new_n230), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(KEYINPUT7), .A3(new_n323), .A4(new_n317), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n319), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(new_n365), .A3(new_n348), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n350), .A2(new_n368), .A3(new_n295), .ZN(new_n369));
  OAI21_X1  g183(.A(G210), .B1(G237), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n350), .A2(new_n368), .A3(new_n295), .A4(new_n370), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n310), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n305), .A2(new_n375), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(G122), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n353), .A2(new_n354), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n220), .B1(new_n378), .B2(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n326), .A2(G122), .A3(new_n327), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(G116), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT88), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(KEYINPUT88), .A3(new_n383), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n203), .A2(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n259), .A2(G143), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G134), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n188), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n380), .A2(new_n220), .A3(new_n382), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n380), .A2(new_n382), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n220), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n390), .B1(new_n389), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n389), .A2(new_n400), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n389), .A2(KEYINPUT87), .A3(new_n400), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n393), .B1(new_n406), .B2(new_n188), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n376), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n394), .A2(new_n395), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n386), .B2(new_n387), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n399), .A2(new_n407), .ZN(new_n412));
  INV_X1    g226(.A(new_n376), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n295), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n397), .A2(new_n408), .A3(new_n376), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n413), .B1(new_n411), .B2(new_n412), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n269), .A2(G952), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(G234), .B2(G237), .ZN(new_n425));
  NAND2_X1  g239(.A1(G234), .A2(G237), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(G902), .A3(G953), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(G898), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(new_n423), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NOR2_X1   g247(.A1(G237), .A2(G953), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G214), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n203), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n434), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT18), .A3(G131), .ZN(new_n440));
  XNOR2_X1  g254(.A(G125), .B(G140), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n201), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT72), .A2(G125), .ZN(new_n443));
  INV_X1    g257(.A(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n442), .B1(new_n447), .B2(new_n201), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n449), .A3(new_n438), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n445), .A2(KEYINPUT16), .A3(new_n446), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT16), .B1(new_n444), .B2(G125), .ZN(new_n453));
  OAI21_X1  g267(.A(G146), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n439), .A2(G131), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n195), .B1(new_n437), .B2(new_n438), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n458), .B2(new_n447), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G146), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n451), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n217), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n456), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(KEYINPUT17), .ZN(new_n468));
  OR3_X1    g282(.A1(new_n452), .A2(G146), .A3(new_n453), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n454), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n464), .B(new_n451), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G475), .A2(G902), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n433), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  AOI211_X1 g289(.A(KEYINPUT20), .B(new_n475), .C1(new_n466), .C2(new_n471), .ZN(new_n476));
  INV_X1    g290(.A(G475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n451), .B1(new_n467), .B2(new_n470), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n465), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n479), .B2(new_n471), .ZN(new_n480));
  OAI22_X1  g294(.A1(new_n474), .A2(new_n476), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n432), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n304), .A2(new_n308), .A3(new_n374), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n336), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n199), .A2(new_n247), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n196), .B(KEYINPUT65), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n190), .A2(G134), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n192), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n260), .A2(new_n261), .B1(G131), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n486), .B1(new_n494), .B2(KEYINPUT30), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n197), .A2(new_n198), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n490), .A2(G131), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n205), .B2(new_n229), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(KEYINPUT66), .A3(new_n491), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n487), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n502), .A2(KEYINPUT67), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT67), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n434), .A2(G210), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT27), .Z(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  OAI211_X1 g324(.A(new_n492), .B(new_n486), .C1(new_n256), .C2(new_n313), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT31), .ZN(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n514), .A2(KEYINPUT28), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n336), .B2(new_n502), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n510), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n506), .A2(new_n521), .A3(new_n510), .A4(new_n511), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(G472), .A2(G902), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT70), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n525), .A2(new_n528), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n506), .A2(new_n531), .A3(new_n519), .A4(new_n511), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n531), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n510), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n511), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n493), .A2(new_n336), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n487), .A2(KEYINPUT71), .A3(new_n486), .A4(new_n492), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n531), .B1(new_n540), .B2(new_n515), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n295), .B(new_n532), .C1(new_n534), .C2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n523), .A2(new_n530), .B1(new_n542), .B2(G472), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n529), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n375), .B1(G234), .B2(new_n295), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n469), .A2(new_n454), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n329), .B2(G128), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n549), .B(new_n550), .C1(G119), .C2(new_n259), .ZN(new_n551));
  XNOR2_X1  g365(.A(G119), .B(G128), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT24), .B(G110), .Z(new_n553));
  AOI22_X1  g367(.A1(new_n551), .A2(G110), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n551), .A2(G110), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n454), .A3(new_n442), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n558), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n295), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(KEYINPUT25), .A3(new_n295), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n546), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n546), .A2(new_n295), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT73), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n570), .B2(new_n562), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n372), .A2(new_n373), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n572), .A2(new_n482), .A3(new_n309), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(KEYINPUT89), .A3(new_n308), .A4(new_n304), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n485), .A2(new_n544), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(G3));
  NAND2_X1  g390(.A1(new_n419), .A2(new_n420), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n419), .A2(KEYINPUT92), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT33), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n419), .B(new_n420), .C1(KEYINPUT92), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(G478), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n416), .A2(new_n295), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n421), .B2(new_n416), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n481), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n372), .A2(KEYINPUT90), .A3(new_n373), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n369), .A2(new_n590), .A3(new_n371), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n309), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n588), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n372), .A2(KEYINPUT90), .A3(new_n373), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n594), .A2(KEYINPUT91), .A3(new_n309), .A4(new_n591), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n593), .A2(new_n431), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n523), .A2(new_n295), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n597), .A2(G472), .B1(new_n526), .B2(new_n523), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n571), .A2(new_n304), .A3(new_n308), .ZN(new_n599));
  AND4_X1   g413(.A1(new_n587), .A2(new_n596), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT34), .B(G104), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NAND2_X1  g416(.A1(new_n418), .A2(new_n423), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n586), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AND4_X1   g419(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n220), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  INV_X1    g423(.A(new_n561), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n558), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n570), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n567), .A2(new_n614), .A3(KEYINPUT94), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT94), .B1(new_n567), .B2(new_n614), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n485), .A2(new_n574), .A3(new_n598), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT37), .B(G110), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G12));
  INV_X1    g435(.A(new_n603), .ZN(new_n622));
  INV_X1    g436(.A(G900), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n425), .B1(new_n428), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n622), .A2(new_n481), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n544), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n304), .A2(new_n308), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n618), .A2(new_n627), .A3(new_n593), .A4(new_n595), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n259), .ZN(G30));
  XOR2_X1   g444(.A(new_n624), .B(KEYINPUT39), .Z(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT40), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n519), .B1(new_n506), .B2(new_n511), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n295), .B1(new_n539), .B2(new_n510), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(KEYINPUT95), .B(G472), .C1(new_n634), .C2(new_n635), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n638), .A2(new_n639), .B1(new_n523), .B2(new_n530), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n640), .A2(new_n529), .A3(KEYINPUT96), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT96), .B1(new_n640), .B2(new_n529), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n572), .B(KEYINPUT38), .Z(new_n644));
  NOR2_X1   g458(.A1(new_n586), .A2(new_n622), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n616), .A2(new_n309), .A3(new_n617), .A4(new_n645), .ZN(new_n646));
  OR4_X1    g460(.A1(new_n633), .A2(new_n643), .A3(new_n644), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G143), .ZN(G45));
  INV_X1    g462(.A(new_n628), .ZN(new_n649));
  INV_X1    g463(.A(new_n624), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n481), .A2(new_n582), .A3(new_n584), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n544), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  INV_X1    g467(.A(new_n571), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n529), .B2(new_n543), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n301), .A2(new_n302), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(G902), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n308), .B(new_n303), .C1(new_n657), .C2(new_n286), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT97), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(new_n596), .A3(new_n659), .A4(new_n587), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  NAND4_X1  g476(.A1(new_n655), .A2(new_n596), .A3(new_n659), .A4(new_n605), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G116), .ZN(G18));
  INV_X1    g478(.A(new_n658), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n593), .A2(new_n665), .A3(new_n595), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(new_n544), .A3(new_n482), .A4(new_n618), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  NAND2_X1  g482(.A1(new_n597), .A2(G472), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n540), .A2(new_n515), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n513), .B(new_n522), .C1(new_n510), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n525), .B(KEYINPUT98), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n669), .A2(new_n571), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n593), .A2(new_n595), .A3(new_n645), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n659), .A4(new_n431), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G122), .ZN(G24));
  AND2_X1   g491(.A1(new_n666), .A2(new_n651), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n597), .A2(G472), .B1(new_n671), .B2(new_n672), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n679), .A2(new_n618), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n679), .B2(new_n618), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  NOR2_X1   g498(.A1(new_n307), .A2(new_n310), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n372), .A2(new_n373), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n268), .A2(new_n687), .A3(new_n274), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n268), .B2(new_n274), .ZN(new_n689));
  OAI211_X1 g503(.A(G469), .B(new_n284), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(G469), .A2(G902), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT100), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n303), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n686), .A2(new_n651), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n523), .A2(new_n530), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n542), .A2(G472), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT32), .B1(new_n523), .B2(new_n526), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n695), .B(new_n571), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n544), .A2(KEYINPUT102), .A3(new_n571), .A4(new_n695), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n700), .B2(new_n703), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT42), .B1(new_n700), .B2(new_n701), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n708), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT104), .B(G131), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G33));
  AND3_X1   g527(.A1(new_n625), .A2(new_n686), .A3(new_n694), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n714), .B(new_n571), .C1(new_n698), .C2(new_n699), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n655), .A2(KEYINPUT105), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  NOR2_X1   g534(.A1(new_n572), .A2(new_n310), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n585), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(KEYINPUT107), .B2(KEYINPUT43), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n724), .B(new_n586), .C1(KEYINPUT107), .C2(new_n723), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n586), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(KEYINPUT106), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n725), .A2(new_n618), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n598), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n722), .B1(new_n732), .B2(KEYINPUT44), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n293), .A2(KEYINPUT45), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n286), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT45), .B(new_n284), .C1(new_n688), .C2(new_n689), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n693), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n303), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n308), .B(new_n631), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n733), .B(new_n744), .C1(KEYINPUT44), .C2(new_n732), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  OAI21_X1  g560(.A(new_n308), .B1(new_n741), .B2(new_n742), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n654), .A2(new_n651), .A3(new_n721), .ZN(new_n752));
  OR3_X1    g566(.A1(new_n751), .A2(new_n544), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  OR2_X1    g568(.A1(new_n681), .A2(new_n682), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n629), .B1(new_n755), .B2(new_n678), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n567), .A2(new_n307), .A3(new_n614), .A4(new_n624), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(new_n694), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n675), .B(new_n759), .C1(new_n641), .C2(new_n642), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n757), .A3(new_n652), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n629), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n683), .A2(new_n762), .A3(new_n760), .A4(new_n652), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n604), .B1(new_n586), .B2(new_n585), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n374), .A2(new_n431), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n599), .A2(new_n598), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n575), .A2(new_n619), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n575), .A2(new_n619), .A3(KEYINPUT109), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n660), .A2(new_n676), .A3(new_n663), .A4(new_n667), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n700), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT103), .B1(new_n778), .B2(KEYINPUT42), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n705), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n709), .A2(KEYINPUT103), .A3(new_n704), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n695), .B1(new_n681), .B2(new_n682), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n721), .A2(new_n586), .A3(new_n622), .A4(new_n650), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n529), .B2(new_n543), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n618), .A2(new_n627), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n717), .A2(new_n718), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n777), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n786), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n766), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n788), .B1(new_n777), .B2(new_n787), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n786), .A2(new_n782), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n791), .A2(new_n711), .A3(KEYINPUT110), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n765), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT111), .B1(new_n800), .B2(KEYINPUT53), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n802));
  NOR2_X1   g616(.A1(new_n777), .A2(new_n787), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n756), .A2(new_n757), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n766), .A2(new_n803), .A3(KEYINPUT53), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n796), .A2(new_n801), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n793), .A2(new_n795), .ZN(new_n807));
  INV_X1    g621(.A(new_n804), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n800), .B1(KEYINPUT53), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n644), .A2(new_n310), .A3(new_n665), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT114), .Z(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(KEYINPUT115), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n725), .A2(new_n425), .A3(new_n730), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n674), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n816), .B(new_n819), .C1(KEYINPUT115), .C2(new_n815), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n665), .A2(new_n721), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n755), .A2(new_n822), .A3(new_n817), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(KEYINPUT115), .B(new_n815), .C1(new_n816), .C2(new_n819), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n643), .A2(new_n571), .A3(new_n425), .A4(new_n822), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n586), .A3(new_n585), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n303), .B1(new_n657), .B2(new_n286), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n751), .B1(new_n308), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n818), .A2(new_n722), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n826), .A2(new_n830), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n830), .A4(new_n836), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n828), .A2(new_n587), .A3(new_n829), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n819), .A2(new_n666), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT117), .Z(new_n843));
  NAND3_X1  g657(.A1(new_n817), .A2(new_n655), .A3(new_n822), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(KEYINPUT48), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n845), .A2(KEYINPUT48), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n424), .B1(new_n844), .B2(new_n846), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n841), .A2(new_n843), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n839), .A2(new_n840), .A3(new_n850), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n812), .A2(new_n851), .B1(G952), .B2(G953), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n654), .A2(new_n728), .A3(new_n307), .A4(new_n310), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n853), .B(new_n644), .C1(KEYINPUT49), .C2(new_n831), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(KEYINPUT49), .B2(new_n831), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n643), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT108), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(G75));
  NAND3_X1  g676(.A1(new_n796), .A2(new_n801), .A3(new_n805), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G210), .A3(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n349), .A2(new_n346), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n325), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n269), .A2(G952), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G51));
  INV_X1    g686(.A(new_n802), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n806), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n863), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n692), .B(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n656), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n863), .A2(G902), .A3(new_n736), .A4(new_n735), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(G54));
  NAND4_X1  g697(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n884));
  INV_X1    g698(.A(new_n472), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n871), .ZN(G60));
  NAND2_X1  g702(.A1(new_n579), .A2(new_n581), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n583), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n889), .A2(new_n875), .A3(new_n877), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n889), .B1(new_n812), .B2(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n871), .A3(new_n893), .ZN(G63));
  NAND2_X1  g708(.A1(G217), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT60), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n612), .B(KEYINPUT122), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n863), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT123), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n863), .A2(new_n900), .A3(new_n896), .A4(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n562), .B1(new_n863), .B2(new_n896), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n871), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n902), .A2(KEYINPUT61), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(G66));
  OAI21_X1  g723(.A(G953), .B1(new_n320), .B2(new_n429), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n791), .B2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n866), .B1(G898), .B2(new_n269), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G69));
  OAI22_X1  g727(.A1(new_n504), .A2(new_n505), .B1(new_n503), .B2(new_n493), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT124), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n460), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n756), .A2(new_n652), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n647), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n655), .A2(new_n721), .A3(new_n767), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(new_n632), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n745), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(new_n753), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n916), .B1(new_n924), .B2(new_n269), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n916), .B1(new_n623), .B2(new_n269), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n744), .A2(new_n655), .A3(new_n675), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n745), .A2(new_n927), .A3(new_n719), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n711), .A2(new_n753), .A3(new_n917), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(new_n269), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n925), .A2(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n931), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G72));
  INV_X1    g749(.A(new_n634), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n506), .A2(new_n519), .A3(new_n511), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n938));
  NAND2_X1  g752(.A1(G472), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n810), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n924), .A2(new_n777), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n936), .B1(new_n944), .B2(new_n941), .ZN(new_n945));
  INV_X1    g759(.A(new_n871), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n929), .B2(new_n791), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n937), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n943), .B(new_n945), .C1(new_n949), .C2(new_n950), .ZN(G57));
endmodule


