//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n210), .B1(new_n211), .B2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n213), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n203), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n217), .B(new_n227), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(KEYINPUT68), .B(G58), .Z(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT8), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(KEYINPUT8), .B2(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n229), .A2(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n228), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n261), .A3(new_n228), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n213), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n257), .A2(new_n264), .B1(new_n201), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n264), .A2(new_n267), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n229), .A2(G1), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(G50), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n276), .B1(new_n277), .B2(new_n274), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n228), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G274), .B1(new_n281), .B2(new_n228), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n282), .A2(new_n287), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT66), .B(G226), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n283), .A2(new_n284), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n283), .A2(new_n293), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n273), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n273), .B(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(G200), .B2(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n299), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n277), .B2(new_n256), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n264), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n267), .A2(new_n203), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n269), .A2(G68), .A3(new_n271), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n274), .A2(new_n275), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n318), .B1(new_n319), .B2(new_n206), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n282), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n290), .B1(G238), .B2(new_n291), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n323), .B2(new_n325), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n317), .B1(new_n329), .B2(G190), .ZN(new_n330));
  INV_X1    g0130(.A(new_n328), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n326), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(G179), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n317), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n269), .A2(G77), .A3(new_n271), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n256), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n264), .B1(new_n277), .B2(new_n267), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n291), .A2(G244), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n289), .B2(new_n288), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n351), .B1(new_n207), .B2(new_n274), .C1(new_n278), .C2(new_n219), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n282), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n343), .B(new_n348), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT69), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(new_n343), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n352), .A2(new_n282), .ZN(new_n360));
  INV_X1    g0160(.A(new_n350), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n359), .A2(KEYINPUT69), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n357), .B(new_n364), .C1(new_n301), .C2(new_n362), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n353), .A2(new_n284), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n366), .B(new_n358), .C1(G169), .C2(new_n353), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n308), .A2(new_n342), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n255), .A2(new_n270), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n269), .B1(new_n267), .B2(new_n255), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n253), .A2(KEYINPUT72), .A3(G68), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT68), .B(G58), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n203), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n231), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n274), .B2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G33), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n386), .A3(KEYINPUT71), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(G68), .C1(KEYINPUT71), .C2(new_n381), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n264), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n274), .A2(new_n380), .A3(G20), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n385), .B2(new_n229), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT16), .B1(new_n379), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n373), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n274), .A2(G226), .A3(G1698), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n396), .B1(new_n319), .B2(new_n220), .C1(new_n320), .C2(new_n279), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n282), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n290), .B1(G232), .B2(new_n291), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G179), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n399), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n405), .B(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n354), .B1(new_n398), .B2(new_n399), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(G190), .B2(new_n400), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n373), .C1(new_n390), .C2(new_n394), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n371), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G116), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n258), .A2(new_n228), .B1(G20), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G283), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n229), .C1(G33), .C2(new_n206), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(KEYINPUT20), .A3(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G1), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G33), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n263), .A2(G116), .A3(new_n266), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n265), .A2(G20), .A3(new_n414), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n286), .A2(G1), .ZN(new_n428));
  AND2_X1   g0228(.A1(KEYINPUT5), .A2(G41), .ZN(new_n429));
  NOR2_X1   g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n289), .ZN(new_n432));
  OR2_X1    g0232(.A1(KEYINPUT5), .A2(G41), .ZN(new_n433));
  NAND2_X1  g0233(.A1(KEYINPUT5), .A2(G41), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n282), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n436), .B2(G270), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n383), .A2(G33), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n439));
  OAI21_X1  g0239(.A(G303), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n382), .A2(new_n384), .A3(G264), .A4(G1698), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n382), .A2(new_n384), .A3(G257), .A4(new_n275), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n282), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n427), .A2(new_n445), .A3(G169), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT21), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(G200), .ZN(new_n449));
  INV_X1    g0249(.A(new_n427), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(G190), .A3(new_n444), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n427), .A2(G179), .A3(new_n444), .A4(new_n437), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n427), .A2(new_n445), .A3(KEYINPUT21), .A4(G169), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n448), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT76), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n454), .A2(new_n453), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(KEYINPUT76), .A3(new_n448), .A4(new_n452), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT74), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n423), .A2(G45), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n289), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G1), .B(G13), .C1(new_n319), .C2(new_n285), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT74), .A3(G274), .A4(new_n428), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(G250), .A3(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n219), .A2(new_n275), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n275), .A2(G244), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n274), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n284), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G169), .B2(new_n473), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT75), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n474), .B(KEYINPUT75), .C1(G169), .C2(new_n473), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n274), .A2(new_n229), .A3(G68), .ZN(new_n479));
  NAND3_X1  g0279(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n229), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G87), .B2(new_n208), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n256), .A2(new_n206), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n479), .B(new_n482), .C1(KEYINPUT19), .C2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n264), .B1(new_n267), .B2(new_n346), .ZN(new_n485));
  INV_X1    g0285(.A(new_n262), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n261), .B1(new_n258), .B2(new_n228), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n266), .B(new_n424), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n346), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n477), .A2(new_n478), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(G87), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n473), .A2(G190), .ZN(new_n496));
  OAI21_X1  g0296(.A(G200), .B1(new_n467), .B2(new_n472), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n220), .A2(KEYINPUT77), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n274), .A2(new_n229), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n274), .A2(KEYINPUT22), .A3(new_n229), .A4(new_n500), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n471), .A2(G20), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT23), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n229), .B2(G107), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n503), .A2(new_n512), .A3(new_n504), .A4(new_n509), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n263), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n266), .A2(G107), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n515), .B(KEYINPUT25), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n207), .B2(new_n488), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n431), .A2(G264), .A3(new_n464), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n221), .A2(G1698), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n382), .A3(new_n384), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT78), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G294), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n382), .A2(new_n384), .A3(G257), .A4(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT78), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n520), .A2(new_n382), .A3(new_n384), .A4(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n519), .B1(new_n527), .B2(new_n282), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n435), .A2(new_n464), .A3(G274), .A4(new_n428), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n301), .A3(new_n529), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n432), .B(new_n519), .C1(new_n527), .C2(new_n282), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G200), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n518), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n529), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n296), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n284), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n514), .C2(new_n517), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n431), .A2(new_n464), .ZN(new_n538));
  INV_X1    g0338(.A(G257), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n529), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n382), .A2(new_n384), .A3(G244), .A4(new_n275), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(KEYINPUT73), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n382), .A2(new_n384), .A3(G250), .A4(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n416), .B(new_n546), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT73), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n284), .B(new_n541), .C1(new_n549), .C2(new_n464), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n251), .A2(G77), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n552), .A2(new_n206), .A3(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(G97), .B(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n555), .B2(new_n229), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n207), .B1(new_n381), .B2(new_n386), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n264), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n267), .A2(new_n206), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n489), .A2(G97), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n542), .A2(new_n543), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT73), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n546), .A2(new_n416), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n564), .A2(new_n544), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n540), .B1(new_n567), .B2(new_n282), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n550), .B(new_n561), .C1(G169), .C2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G190), .B(new_n541), .C1(new_n549), .C2(new_n464), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n559), .B1(new_n488), .B2(new_n206), .ZN(new_n571));
  OAI21_X1  g0371(.A(G107), .B1(new_n391), .B2(new_n392), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n554), .A2(new_n552), .ZN(new_n573));
  INV_X1    g0373(.A(new_n553), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G20), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n551), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n571), .B1(new_n577), .B2(new_n264), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n570), .B(new_n578), .C1(new_n354), .C2(new_n568), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n533), .A2(new_n537), .A3(new_n569), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n499), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n413), .A2(new_n460), .A3(new_n581), .ZN(G372));
  NAND2_X1  g0382(.A1(new_n341), .A2(new_n317), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n335), .B2(new_n367), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n411), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n407), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n305), .A2(new_n307), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n298), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n585), .A2(new_n407), .B1(new_n305), .B2(new_n307), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n299), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n413), .ZN(new_n594));
  INV_X1    g0394(.A(new_n467), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n470), .A2(new_n471), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n282), .ZN(new_n598));
  AOI211_X1 g0398(.A(KEYINPUT79), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(new_n296), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n492), .A2(new_n474), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n537), .A2(new_n448), .A3(new_n458), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n537), .A2(KEYINPUT82), .A3(new_n458), .A4(new_n448), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n533), .A2(new_n569), .A3(new_n579), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(G200), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT80), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n485), .A2(new_n612), .A3(new_n494), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n485), .B2(new_n494), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(KEYINPUT81), .B1(G190), .B2(new_n473), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT81), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n611), .B(new_n617), .C1(new_n613), .C2(new_n614), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n603), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n604), .B1(new_n610), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g0421(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n499), .A2(new_n569), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n615), .A2(KEYINPUT81), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n496), .A3(new_n618), .ZN(new_n626));
  INV_X1    g0426(.A(new_n569), .ZN(new_n627));
  INV_X1    g0427(.A(new_n603), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n593), .B1(new_n594), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT86), .ZN(G369));
  NAND2_X1  g0433(.A1(new_n458), .A2(new_n448), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n265), .A2(new_n229), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n450), .A2(new_n641), .ZN(new_n642));
  MUX2_X1   g0442(.A(new_n460), .B(new_n634), .S(new_n642), .Z(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G330), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n533), .B(new_n537), .C1(new_n518), .C2(new_n641), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n537), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n640), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n644), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n640), .B1(new_n458), .B2(new_n448), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n641), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n652), .A2(new_n656), .ZN(G399));
  NAND2_X1  g0457(.A1(new_n215), .A2(new_n285), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT88), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n220), .A2(new_n206), .A3(new_n207), .A4(new_n414), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n659), .A2(new_n423), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n233), .B2(new_n659), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT28), .Z(new_n663));
  NOR3_X1   g0463(.A1(new_n631), .A2(KEYINPUT29), .A3(new_n640), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT29), .ZN(new_n665));
  INV_X1    g0465(.A(new_n604), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n609), .A2(new_n605), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n668), .B2(new_n619), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n619), .A2(KEYINPUT26), .A3(new_n627), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n622), .B1(new_n499), .B2(new_n569), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n665), .B1(new_n673), .B2(new_n641), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n547), .A2(new_n548), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n464), .B1(new_n677), .B2(new_n544), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n437), .A2(G179), .A3(new_n444), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n678), .A2(new_n679), .A3(new_n540), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n528), .A2(new_n473), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT89), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n528), .A2(new_n473), .A3(KEYINPUT89), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n443), .A2(new_n282), .ZN(new_n686));
  INV_X1    g0486(.A(G270), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n529), .B1(new_n538), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n284), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n531), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n568), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n600), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT90), .B(new_n595), .C1(new_n598), .C2(new_n599), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n690), .A2(new_n691), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n686), .A2(new_n284), .A3(new_n688), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n568), .A2(new_n697), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n528), .A2(new_n473), .A3(KEYINPUT89), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT89), .B1(new_n528), .B2(new_n473), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT91), .B1(new_n701), .B2(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n680), .A2(new_n684), .A3(new_n683), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n696), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT31), .B1(new_n707), .B2(new_n640), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n705), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n709), .B(new_n641), .C1(new_n696), .C2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n676), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n696), .A2(new_n710), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n685), .A2(new_n695), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n641), .B1(new_n717), .B2(new_n706), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT92), .B(new_n714), .C1(new_n718), .C2(KEYINPUT31), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n533), .A2(new_n537), .A3(new_n569), .A4(new_n579), .ZN(new_n720));
  INV_X1    g0520(.A(new_n498), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n475), .A2(new_n476), .B1(new_n491), .B2(new_n485), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n478), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n460), .A2(new_n720), .A3(new_n723), .A4(new_n641), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT93), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n460), .A4(new_n641), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n712), .A2(new_n719), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n675), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n663), .B1(new_n732), .B2(G1), .ZN(G364));
  XOR2_X1   g0533(.A(new_n644), .B(KEYINPUT94), .Z(new_n734));
  NOR2_X1   g0534(.A1(new_n213), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n423), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n659), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n734), .B(new_n739), .C1(G330), .C2(new_n643), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n228), .B1(G20), .B2(new_n296), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n249), .A2(G45), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT95), .Z(new_n748));
  INV_X1    g0548(.A(new_n215), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n274), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n748), .B(new_n750), .C1(G45), .C2(new_n232), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G355), .A2(new_n274), .ZN(new_n752));
  MUX2_X1   g0552(.A(G116), .B(new_n752), .S(new_n215), .Z(new_n753));
  AOI21_X1  g0553(.A(new_n746), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G20), .A2(G179), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G190), .A3(new_n354), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G322), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G326), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n229), .A2(G179), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(new_n301), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G329), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n767), .A2(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n765), .B1(KEYINPUT98), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(KEYINPUT98), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n756), .A2(new_n769), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n301), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n229), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n385), .B1(new_n778), .B2(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n354), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n756), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n777), .B(new_n783), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n763), .A2(new_n774), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n778), .A2(new_n220), .ZN(new_n790));
  INV_X1    g0590(.A(new_n781), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G97), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  OAI21_X1  g0593(.A(KEYINPUT32), .B1(new_n770), .B2(new_n793), .ZN(new_n794));
  OR3_X1    g0594(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n793), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n764), .B2(G50), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n274), .B1(new_n207), .B2(new_n767), .C1(new_n775), .C2(new_n277), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G68), .B2(new_n787), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(new_n376), .C2(new_n761), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n739), .B(new_n754), .C1(new_n744), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n743), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n643), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n740), .A2(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n358), .A2(new_n640), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n355), .A2(new_n356), .B1(new_n301), .B2(new_n362), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT69), .B1(new_n359), .B2(new_n363), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n367), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT100), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT100), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n365), .A2(new_n811), .A3(new_n367), .A4(new_n806), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n367), .A2(new_n641), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n631), .B2(new_n640), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n812), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n641), .B(new_n816), .C1(new_n621), .C2(new_n630), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n738), .B1(new_n818), .B2(new_n730), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n730), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n744), .A2(new_n741), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n738), .B1(G77), .B2(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n414), .A2(new_n775), .B1(new_n786), .B2(new_n768), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n385), .B1(new_n770), .B2(new_n776), .C1(new_n781), .C2(new_n206), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n220), .A2(new_n767), .B1(new_n778), .B2(new_n207), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n764), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n779), .B2(new_n828), .C1(new_n761), .C2(new_n782), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT99), .Z(new_n830));
  INV_X1    g0630(.A(new_n775), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G150), .A2(new_n787), .B1(new_n831), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n828), .C1(new_n761), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n274), .B1(new_n770), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n781), .A2(new_n376), .B1(new_n767), .B2(new_n203), .ZN(new_n840));
  INV_X1    g0640(.A(new_n778), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n840), .C1(G50), .C2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n835), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(KEYINPUT34), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n830), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n823), .B1(new_n845), .B2(new_n744), .ZN(new_n846));
  INV_X1    g0646(.A(new_n814), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n742), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n820), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n230), .A2(G116), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n575), .B2(KEYINPUT35), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(KEYINPUT35), .B2(new_n575), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT36), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n374), .A2(new_n377), .A3(G77), .A4(new_n233), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(G50), .B2(new_n203), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(G1), .A3(new_n213), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT101), .Z(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n379), .B2(new_n388), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n373), .B1(new_n390), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n638), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT103), .B(new_n373), .C1(new_n390), .C2(new_n860), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT104), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n863), .A2(KEYINPUT104), .A3(new_n864), .A4(new_n865), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n863), .A2(new_n404), .A3(new_n865), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n868), .A2(new_n410), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n395), .A2(new_n864), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n405), .A2(new_n872), .A3(new_n410), .A4(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n405), .A2(new_n410), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n873), .A4(new_n872), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n871), .A2(KEYINPUT37), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n407), .A2(new_n411), .B1(new_n868), .B2(new_n869), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n876), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n872), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n872), .B1(new_n407), .B2(new_n411), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n583), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n341), .A2(KEYINPUT102), .A3(new_n317), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n330), .A2(new_n333), .B1(new_n317), .B2(new_n640), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n317), .B(new_n640), .C1(new_n335), .C2(new_n341), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n814), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n707), .A2(new_n640), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(new_n709), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n726), .A2(new_n727), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT40), .B1(new_n890), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(KEYINPUT107), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n883), .ZN(new_n905));
  INV_X1    g0705(.A(new_n881), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(KEYINPUT40), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n903), .B(new_n909), .C1(new_n901), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n899), .A2(new_n900), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n913), .A2(new_n413), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(new_n413), .B2(new_n914), .ZN(new_n916));
  INV_X1    g0716(.A(G330), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n882), .B2(new_n889), .ZN(new_n920));
  INV_X1    g0720(.A(new_n893), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT102), .B1(new_n341), .B2(new_n317), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n641), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT106), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n920), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n407), .A2(new_n864), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n895), .A2(new_n896), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n367), .A2(new_n640), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n817), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n927), .B1(new_n909), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n413), .B1(new_n664), .B2(new_n674), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n593), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n918), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n918), .A2(new_n937), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT108), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n938), .B1(new_n423), .B2(new_n735), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n939), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n859), .B1(new_n941), .B2(new_n943), .ZN(G367));
  NOR2_X1   g0744(.A1(new_n778), .A2(new_n414), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n786), .A2(new_n782), .B1(new_n945), .B2(KEYINPUT46), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT46), .ZN(new_n947));
  INV_X1    g0747(.A(new_n767), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(G97), .ZN(new_n949));
  INV_X1    g0749(.A(new_n770), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n274), .B1(new_n950), .B2(G317), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n946), .B(new_n952), .C1(G311), .C2(new_n764), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n775), .A2(new_n768), .B1(new_n207), .B2(new_n781), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT110), .Z(new_n955));
  OAI211_X1 g0755(.A(new_n953), .B(new_n955), .C1(new_n779), .C2(new_n761), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n201), .A2(new_n775), .B1(new_n786), .B2(new_n793), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n274), .B1(new_n770), .B2(new_n833), .C1(new_n376), .C2(new_n778), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n781), .A2(new_n203), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n767), .A2(new_n277), .ZN(new_n960));
  NOR4_X1   g0760(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(G150), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n961), .B1(new_n834), .B2(new_n828), .C1(new_n962), .C2(new_n761), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n744), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n750), .A2(new_n242), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n745), .C1(new_n215), .C2(new_n346), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n738), .A3(new_n968), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n613), .A2(new_n614), .A3(new_n641), .ZN(new_n970));
  MUX2_X1   g0770(.A(new_n620), .B(new_n604), .S(new_n970), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n969), .B1(new_n743), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n627), .A2(new_n640), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n569), .B(new_n579), .C1(new_n578), .C2(new_n641), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n656), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT44), .Z(new_n978));
  NAND3_X1  g0778(.A1(new_n654), .A2(new_n655), .A3(new_n975), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n981), .A2(new_n982), .B1(new_n652), .B2(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n652), .A2(KEYINPUT109), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n978), .B(new_n983), .C1(KEYINPUT109), .C2(new_n652), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n649), .A2(new_n651), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n654), .B1(new_n989), .B2(new_n653), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n644), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n734), .B2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n731), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n659), .B(KEYINPUT41), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n736), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n971), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n654), .A2(new_n976), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT42), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n974), .A2(new_n537), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n640), .B1(new_n1000), .B2(new_n569), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n998), .B2(KEYINPUT42), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n997), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n971), .A2(new_n996), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n652), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n976), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1008), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n972), .B1(new_n995), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(G387));
  AND3_X1   g0813(.A1(new_n239), .A2(G45), .A3(new_n385), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n344), .A2(new_n201), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1017));
  AOI21_X1  g0817(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n660), .B1(new_n1019), .B2(new_n385), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n215), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n746), .B1(G107), .B2(new_n749), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n739), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n989), .B2(new_n803), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n761), .A2(new_n201), .B1(new_n346), .B2(new_n781), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT111), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n385), .B1(new_n950), .B2(G150), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n949), .C1(new_n277), .C2(new_n778), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n255), .A2(new_n786), .B1(new_n203), .B2(new_n775), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G159), .C2(new_n764), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n274), .B1(new_n950), .B2(G326), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G303), .A2(new_n831), .B1(new_n787), .B2(G311), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT112), .B(G322), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n828), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G317), .B2(new_n762), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT113), .Z(new_n1037));
  INV_X1    g0837(.A(KEYINPUT48), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n791), .A2(G283), .B1(new_n841), .B2(G294), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1032), .B1(new_n414), .B2(new_n767), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1031), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1024), .B1(new_n1046), .B2(new_n744), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n737), .B2(new_n992), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n732), .A2(new_n992), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n659), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n732), .A2(new_n992), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  AND2_X1   g0852(.A1(new_n732), .A2(new_n992), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n988), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(new_n986), .A3(new_n987), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n659), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n976), .A2(new_n743), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n745), .B1(new_n206), .B2(new_n215), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n246), .B2(new_n750), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n762), .A2(G311), .B1(G317), .B2(new_n764), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n385), .B1(new_n770), .B2(new_n1034), .C1(new_n207), .C2(new_n767), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n781), .A2(new_n414), .B1(new_n778), .B2(new_n768), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n782), .B2(new_n775), .C1(new_n779), .C2(new_n786), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n761), .A2(new_n793), .B1(new_n962), .B2(new_n828), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  AOI22_X1  g0868(.A1(G50), .A2(new_n787), .B1(new_n831), .B2(new_n344), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n274), .B1(new_n770), .B2(new_n834), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G87), .B2(new_n948), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n791), .A2(G77), .B1(new_n841), .B2(G68), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1062), .A2(new_n1066), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n739), .B(new_n1059), .C1(new_n1074), .C2(new_n744), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n988), .A2(new_n737), .B1(new_n1057), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1056), .A2(new_n1076), .ZN(G390));
  NAND3_X1  g0877(.A1(new_n914), .A2(G330), .A3(new_n897), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n924), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n817), .A2(new_n931), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n928), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n920), .A2(new_n925), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n673), .A2(new_n641), .A3(new_n816), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n929), .B1(new_n1084), .B2(new_n931), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n890), .A2(new_n924), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1082), .A2(new_n1080), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n878), .A2(new_n876), .B1(new_n884), .B2(KEYINPUT37), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n880), .B1(new_n1090), .B2(new_n887), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT39), .B1(new_n907), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1088), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n729), .A2(G330), .A3(new_n897), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT115), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n729), .A2(KEYINPUT115), .A3(new_n897), .A4(G330), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1084), .A2(new_n931), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n928), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n1080), .C1(new_n882), .C2(new_n889), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1087), .A2(new_n1102), .A3(new_n737), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n741), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n761), .A2(new_n414), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G97), .A2(new_n831), .B1(new_n787), .B2(G107), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n274), .B(new_n790), .C1(G294), .C2(new_n950), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n764), .A2(G283), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n791), .A2(G77), .B1(new_n948), .B2(G68), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n761), .A2(new_n838), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n274), .B1(new_n770), .B2(new_n1112), .C1(new_n201), .C2(new_n767), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G159), .B2(new_n791), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  NOR2_X1   g0915(.A1(new_n778), .A2(new_n962), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n831), .A2(new_n1115), .B1(new_n1117), .B2(KEYINPUT53), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT53), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n787), .A2(G137), .B1(new_n1119), .B2(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n764), .A2(G128), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1114), .A2(new_n1118), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1105), .A2(new_n1110), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n744), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n255), .A2(new_n821), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1104), .A2(new_n738), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1103), .A2(KEYINPUT117), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT117), .B1(new_n1103), .B2(new_n1126), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1103), .A2(new_n1126), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT118), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1127), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1087), .A2(new_n1102), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n729), .A2(G330), .A3(new_n847), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n929), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1078), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1081), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n847), .C1(new_n899), .C2(new_n900), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1099), .B1(new_n1141), .B2(new_n929), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1098), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n914), .A2(G330), .A3(new_n413), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n935), .A2(new_n593), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT116), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT116), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1149), .B(new_n1146), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1136), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1081), .A2(new_n1139), .B1(new_n1098), .B2(new_n1142), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1149), .B1(new_n1152), .B2(new_n1146), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1087), .A2(new_n1102), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1144), .A2(KEYINPUT116), .A3(new_n1147), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n659), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1130), .A2(new_n1135), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(G378));
  NAND2_X1  g0959(.A1(new_n273), .A2(new_n864), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n308), .B(new_n1160), .Z(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n934), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n926), .A2(new_n933), .A3(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n917), .B1(new_n902), .B2(new_n912), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1168), .A3(new_n1166), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1164), .A2(new_n741), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n791), .A2(G150), .B1(new_n841), .B2(new_n1115), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n775), .B2(new_n833), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G132), .B2(new_n787), .ZN(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1176), .B1(new_n1112), .B2(new_n828), .C1(new_n1177), .C2(new_n761), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT119), .Z(new_n1179));
  AND2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(G33), .A2(G41), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT120), .B(G124), .Z(new_n1183));
  OAI221_X1 g0983(.A(new_n1182), .B1(new_n767), .B2(new_n793), .C1(new_n770), .C2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n206), .A2(new_n786), .B1(new_n775), .B2(new_n346), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n274), .A2(G41), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n768), .B2(new_n770), .C1(new_n203), .C2(new_n781), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n778), .A2(new_n277), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n767), .A2(new_n376), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n207), .B2(new_n761), .C1(new_n414), .C2(new_n828), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1187), .A2(G50), .A3(new_n1182), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n744), .B1(new_n1185), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT121), .Z(new_n1199));
  AOI211_X1 g0999(.A(new_n739), .B(new_n1199), .C1(new_n201), .C2(new_n821), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1172), .A2(new_n737), .B1(new_n1173), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1151), .A2(new_n1147), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1172), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1146), .B1(new_n1204), .B2(new_n1136), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1165), .A2(new_n1168), .A3(new_n1166), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1168), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n659), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1201), .B1(new_n1203), .B2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n929), .A2(new_n741), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n738), .B1(G68), .B2(new_n822), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n761), .A2(new_n768), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G107), .A2(new_n831), .B1(new_n787), .B2(G116), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n274), .B(new_n960), .C1(G303), .C2(new_n950), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n764), .A2(G294), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n791), .A2(new_n490), .B1(new_n841), .B2(G97), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n761), .A2(new_n833), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G150), .A2(new_n831), .B1(new_n787), .B2(new_n1115), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n764), .A2(G132), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n274), .B1(new_n770), .B2(new_n1177), .C1(new_n376), .C2(new_n767), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n791), .A2(G50), .B1(new_n841), .B2(G159), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1213), .A2(new_n1218), .B1(new_n1219), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1212), .B1(new_n1226), .B2(new_n744), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1144), .A2(new_n737), .B1(new_n1211), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1152), .A2(new_n1146), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n994), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1204), .B2(new_n1231), .ZN(G381));
  NAND2_X1  g1032(.A1(new_n1133), .A2(new_n1127), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1012), .A2(new_n849), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G375), .A2(new_n1235), .A3(new_n1238), .A4(G381), .ZN(G407));
  NAND2_X1  g1039(.A1(new_n639), .A2(G213), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(G375), .A2(new_n1235), .A3(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT122), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1043(.A(new_n1228), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n659), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1153), .A2(new_n1155), .A3(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1229), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(KEYINPUT123), .A3(new_n1229), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n849), .B(new_n1244), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1246), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1251), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G384), .B1(new_n1255), .B2(new_n1228), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1154), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1172), .B(new_n1230), .C1(new_n1258), .C2(new_n1146), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1201), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1234), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(G375), .B2(new_n1158), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(new_n1262), .A3(new_n1240), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1240), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1247), .A2(KEYINPUT123), .A3(new_n1229), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT123), .B1(new_n1247), .B2(new_n1229), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1246), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n849), .B1(new_n1268), .B2(new_n1244), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1255), .A2(G384), .A3(new_n1228), .ZN(new_n1270));
  INV_X1    g1070(.A(G2897), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1240), .A2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1265), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1257), .A2(new_n1262), .A3(new_n1277), .A4(new_n1240), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1264), .A2(new_n1275), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(new_n1236), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1012), .A2(G390), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT125), .B1(new_n1012), .B2(G390), .ZN(new_n1283));
  XOR2_X1   g1083(.A(G393), .B(G396), .Z(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1280), .A2(new_n1283), .A3(new_n1281), .A4(new_n1284), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1252), .A2(new_n1256), .B1(new_n1271), .B2(new_n1240), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(KEYINPUT124), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1291), .A2(new_n1265), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1263), .A2(KEYINPUT63), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1257), .A2(new_n1262), .A3(new_n1297), .A4(new_n1240), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT126), .B1(new_n1288), .B2(KEYINPUT61), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1286), .A2(new_n1301), .A3(new_n1276), .A4(new_n1287), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1295), .A2(new_n1299), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1289), .A2(new_n1304), .ZN(G405));
  XNOR2_X1  g1105(.A(new_n1288), .B(new_n1257), .ZN(new_n1306));
  AND2_X1   g1106(.A1(G375), .A2(new_n1234), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT127), .B1(G375), .B2(new_n1158), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1307), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1306), .B(new_n1311), .ZN(G402));
endmodule


