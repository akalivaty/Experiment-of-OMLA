//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973;
  OR2_X1    g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT76), .ZN(new_n206));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT77), .B(G162gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n203), .B1(new_n212), .B2(G155gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n202), .B(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n211), .B(KEYINPUT78), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(G211gat), .A2(G218gat), .ZN(new_n219));
  INV_X1    g018(.A(G211gat), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G197gat), .A2(G204gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G197gat), .A2(G204gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n219), .B(new_n222), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n219), .ZN(new_n228));
  XNOR2_X1  g027(.A(G197gat), .B(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n226), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT29), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n217), .B(new_n218), .C1(KEYINPUT3), .C2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n211), .B(new_n234), .C1(new_n213), .C2(new_n214), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n227), .A2(new_n231), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(G228gat), .A3(new_n240), .A4(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n234), .B1(new_n232), .B2(new_n244), .ZN(new_n245));
  AOI211_X1 g044(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n227), .C2(new_n231), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n215), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n237), .A2(KEYINPUT83), .A3(new_n239), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n250));
  NAND2_X1  g049(.A1(G228gat), .A2(G233gat), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n241), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G22gat), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n256), .B(new_n241), .C1(new_n252), .C2(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G78gat), .B(G106gat), .ZN(new_n259));
  INV_X1    g058(.A(G50gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n263));
  INV_X1    g062(.A(new_n261), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n255), .A2(new_n264), .A3(new_n257), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n263), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n255), .A2(new_n264), .A3(new_n257), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n255), .B2(new_n257), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G227gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G127gat), .B(G134gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G120gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G113gat), .ZN(new_n283));
  INV_X1    g082(.A(G113gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G120gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT68), .A4(new_n279), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n281), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT69), .B1(new_n281), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT27), .B(G183gat), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT28), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT28), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  OAI221_X1 g105(.A(new_n292), .B1(new_n296), .B2(new_n300), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n301), .A2(new_n302), .A3(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(new_n295), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n298), .B2(KEYINPUT23), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT67), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n310), .A2(new_n321), .A3(new_n311), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n315), .A2(G169gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n294), .A2(KEYINPUT64), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G176gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n316), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT65), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(new_n317), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT25), .B1(new_n295), .B2(new_n315), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n297), .B1(new_n298), .B2(KEYINPUT23), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT66), .B(G190gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n310), .B(new_n311), .C1(new_n334), .C2(G183gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n329), .B1(new_n328), .B2(new_n317), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n291), .B(new_n307), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n328), .A2(new_n317), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT65), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(new_n330), .A3(new_n320), .A4(new_n337), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n291), .B1(new_n344), .B2(new_n307), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n276), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT33), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n273), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  INV_X1    g148(.A(new_n276), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n307), .B1(new_n338), .B2(new_n339), .ZN(new_n351));
  INV_X1    g150(.A(new_n291), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n353), .B2(new_n340), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT32), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n346), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n348), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n350), .A3(new_n340), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n346), .B(KEYINPUT32), .C1(new_n347), .C2(new_n273), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n358), .B2(new_n363), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n359), .A2(new_n360), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT34), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n358), .A2(new_n363), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n361), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n372), .B2(new_n364), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n266), .B(new_n270), .C1(new_n370), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n351), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n344), .B2(new_n307), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n239), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n377), .B(new_n238), .C1(new_n378), .C2(new_n376), .ZN(new_n381));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  NAND4_X1  g183(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT30), .A4(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n380), .A2(new_n381), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n384), .B(KEYINPUT72), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT73), .B(new_n390), .C1(new_n380), .C2(new_n381), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n386), .B(new_n387), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n392), .A2(new_n393), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(KEYINPUT75), .A3(new_n386), .A4(new_n387), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n217), .A2(KEYINPUT3), .A3(new_n218), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n281), .A2(new_n288), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n235), .ZN(new_n401));
  INV_X1    g200(.A(new_n215), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n291), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n215), .A2(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n401), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n217), .A2(new_n218), .A3(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n406), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n412), .B2(new_n405), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n215), .A2(new_n400), .A3(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(new_n290), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n281), .A2(new_n288), .A3(KEYINPUT69), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n402), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n415), .B1(new_n418), .B2(new_n407), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n405), .A2(KEYINPUT5), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n401), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n429), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n414), .A2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(new_n427), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n384), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n389), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT30), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n396), .A2(new_n398), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT35), .B1(new_n374), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n270), .A2(new_n266), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n394), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n427), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n434), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n430), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT35), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n438), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n444), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n369), .B1(new_n365), .B2(new_n366), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n372), .A2(new_n364), .A3(new_n368), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n443), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT36), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n404), .B1(new_n419), .B2(new_n401), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT39), .B1(new_n412), .B2(new_n405), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT85), .B(KEYINPUT39), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n427), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n462), .B2(new_n464), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n446), .A2(new_n447), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n394), .B2(new_n438), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n389), .A2(KEYINPUT37), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n380), .A2(new_n381), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n436), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT38), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n390), .A2(KEYINPUT38), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n389), .B2(KEYINPUT37), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n437), .B1(new_n478), .B2(new_n474), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n479), .A3(new_n448), .A4(new_n449), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n471), .A2(new_n270), .A3(new_n266), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n455), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n458), .A2(new_n459), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n457), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G232gat), .A2(G233gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT93), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT41), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT94), .Z(new_n490));
  XNOR2_X1  g289(.A(G134gat), .B(G162gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  INV_X1    g295(.A(G43gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(G50gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n260), .A2(G43gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n496), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n499), .A3(KEYINPUT15), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  INV_X1    g304(.A(G29gat), .ZN(new_n506));
  INV_X1    g305(.A(G36gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G29gat), .A2(G36gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT89), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n503), .A2(new_n504), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n504), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n494), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n512), .A2(new_n504), .A3(new_n510), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n524), .A2(new_n503), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT95), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n531), .A2(G85gat), .A3(G92gat), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G99gat), .B(G106gat), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(G85gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n534), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n536), .B1(new_n534), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n522), .B2(new_n521), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n543), .A2(new_n521), .B1(KEYINPUT41), .B2(new_n488), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n547), .B1(new_n545), .B2(new_n548), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n545), .A2(new_n548), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n546), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n556), .B2(new_n549), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n493), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT98), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT98), .B(new_n493), .C1(new_n554), .C2(new_n557), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n552), .B1(new_n550), .B2(new_n553), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(new_n551), .A3(new_n549), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n492), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT99), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n492), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n560), .A2(new_n561), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n572), .B(new_n571), .C1(new_n569), .C2(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G127gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G15gat), .B(G22gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT16), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(G1gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(G1gat), .B2(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G8gat), .ZN(new_n589));
  INV_X1    g388(.A(G8gat), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n587), .B(new_n590), .C1(G1gat), .C2(new_n585), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n579), .B2(new_n578), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n584), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G155gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n594), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n568), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G197gat), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT11), .B(G169gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n591), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n522), .B2(new_n521), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n527), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n521), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n608), .A2(KEYINPUT18), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n609), .B(KEYINPUT13), .Z(new_n612));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n613), .A3(new_n525), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n610), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n592), .B2(new_n525), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n527), .A2(new_n607), .B1(new_n606), .B2(new_n521), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT18), .B1(new_n619), .B2(new_n609), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n605), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n605), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n611), .A4(new_n617), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(KEYINPUT92), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT92), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n628), .B(new_n605), .C1(new_n618), .C2(new_n620), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n578), .B1(new_n541), .B2(new_n542), .ZN(new_n631));
  INV_X1    g430(.A(new_n533), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n531), .A2(new_n532), .B1(G85gat), .B2(G92gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n540), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n535), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n576), .A2(new_n577), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n534), .A2(new_n536), .A3(new_n540), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n631), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n543), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n631), .A2(new_n638), .ZN(new_n645));
  INV_X1    g444(.A(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT100), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n644), .A2(new_n647), .A3(new_n654), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n652), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n600), .A2(new_n630), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n485), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n435), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n435), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g466(.A1(new_n444), .A2(new_n451), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AND3_X1   g468(.A1(new_n660), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n590), .B1(new_n660), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n670), .ZN(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n660), .A2(new_n674), .A3(new_n455), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n483), .A2(new_n459), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n660), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n442), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n560), .A2(new_n561), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n565), .A2(new_n567), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n485), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n568), .B1(new_n457), .B2(new_n484), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n599), .A2(new_n630), .A3(new_n658), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n665), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n506), .B1(new_n693), .B2(KEYINPUT104), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT104), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n692), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n664), .A2(G29gat), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n696), .A2(KEYINPUT103), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n696), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n695), .A2(new_n702), .ZN(G1328gat));
  NAND3_X1  g502(.A1(new_n691), .A2(new_n668), .A3(new_n692), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n507), .B1(new_n704), .B2(KEYINPUT105), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT105), .B2(new_n704), .ZN(new_n706));
  INV_X1    g505(.A(new_n668), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n696), .A2(G36gat), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT46), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n691), .A2(new_n676), .A3(new_n692), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  INV_X1    g512(.A(new_n696), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n497), .A3(new_n455), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n712), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1330gat));
  NAND3_X1  g517(.A1(new_n691), .A2(new_n442), .A3(new_n692), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G50gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n442), .A2(new_n260), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n714), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n720), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1331gat));
  AND2_X1   g526(.A1(new_n627), .A2(new_n629), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n600), .A2(new_n728), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n485), .A2(new_n658), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n664), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n662), .A2(KEYINPUT108), .A3(new_n663), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n738));
  INV_X1    g537(.A(G64gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n730), .B(new_n668), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT109), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n730), .A2(new_n744), .A3(new_n455), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n730), .A2(new_n676), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n744), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n442), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT110), .B(G78gat), .Z(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1335gat));
  INV_X1    g550(.A(new_n658), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n728), .A2(new_n599), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n691), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n664), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n728), .A2(new_n599), .ZN(new_n756));
  AND4_X1   g555(.A1(KEYINPUT51), .A2(new_n485), .A3(new_n685), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n689), .B2(new_n756), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(new_n538), .A3(new_n665), .A4(new_n658), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(G1336gat));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n707), .A2(G92gat), .A3(new_n752), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n688), .A2(new_n690), .A3(new_n668), .A4(new_n753), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n766), .B(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(new_n676), .ZN(new_n771));
  OAI21_X1  g570(.A(G99gat), .B1(new_n754), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n455), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(G99gat), .A3(new_n752), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(G1338gat));
  NAND4_X1  g575(.A1(new_n688), .A2(new_n690), .A3(new_n442), .A4(new_n753), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n443), .A2(G106gat), .A3(new_n752), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n757), .B2(new_n758), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT112), .B(new_n780), .C1(new_n757), .C2(new_n758), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n778), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n786), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n786), .B2(KEYINPUT53), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(G1339gat));
  NAND4_X1  g588(.A1(new_n568), .A2(new_n599), .A3(new_n630), .A4(new_n752), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT114), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT117), .B1(new_n619), .B2(new_n609), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n615), .A2(new_n616), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n612), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n619), .A2(KEYINPUT117), .A3(new_n609), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n604), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(new_n626), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n646), .B1(new_n640), .B2(new_n641), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI211_X1 g600(.A(KEYINPUT54), .B(new_n646), .C1(new_n640), .C2(new_n641), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n802), .B2(new_n651), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n800), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(new_n652), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n801), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n656), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(new_n801), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n804), .B2(new_n652), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT115), .B(new_n651), .C1(new_n799), .C2(new_n800), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n809), .B(KEYINPUT55), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT116), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n656), .A4(new_n812), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n685), .A2(new_n797), .A3(new_n814), .A4(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n728), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n797), .A2(new_n658), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n685), .B1(new_n824), .B2(KEYINPUT118), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n821), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n791), .B1(new_n828), .B2(new_n599), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n734), .ZN(new_n831));
  INV_X1    g630(.A(new_n374), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n668), .ZN(new_n834));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n728), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n664), .A2(new_n668), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n829), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n630), .A2(new_n284), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(G1340gat));
  AOI21_X1  g638(.A(new_n282), .B1(new_n837), .B2(new_n658), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT119), .Z(new_n841));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n282), .A3(new_n658), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1341gat));
  NAND3_X1  g642(.A1(new_n834), .A2(new_n583), .A3(new_n599), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n837), .A2(new_n599), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n583), .B2(new_n846), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n707), .A2(new_n685), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(G134gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n832), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n837), .A2(new_n685), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n850), .A2(KEYINPUT56), .B1(new_n851), .B2(G134gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n850), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(G1343gat));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n829), .A2(new_n858), .A3(new_n735), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n676), .A2(new_n443), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n858), .B1(new_n829), .B2(new_n735), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n861), .A2(new_n862), .A3(new_n668), .A4(new_n630), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n771), .A2(new_n836), .ZN(new_n864));
  INV_X1    g663(.A(new_n791), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n817), .A2(new_n656), .A3(new_n812), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(new_n630), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n685), .B1(new_n823), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n599), .B1(new_n869), .B2(new_n820), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n442), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n864), .B1(new_n871), .B2(KEYINPUT57), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n829), .A2(new_n873), .A3(new_n442), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n728), .A2(G141gat), .ZN(new_n876));
  OAI22_X1  g675(.A1(new_n863), .A2(G141gat), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI221_X1 g678(.A(KEYINPUT58), .B1(new_n875), .B2(new_n876), .C1(new_n863), .C2(G141gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1344gat));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n862), .ZN(new_n882));
  INV_X1    g681(.A(G148gat), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n707), .A4(new_n658), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n873), .B1(new_n829), .B2(new_n442), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n442), .A2(new_n873), .ZN(new_n887));
  INV_X1    g686(.A(new_n599), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n685), .A2(new_n797), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n866), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n890), .B2(new_n868), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n891), .B2(new_n790), .ZN(new_n892));
  NOR4_X1   g691(.A1(new_n886), .A2(new_n752), .A3(new_n864), .A4(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n883), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n886), .ZN(new_n896));
  INV_X1    g695(.A(new_n864), .ZN(new_n897));
  INV_X1    g696(.A(new_n892), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n896), .A2(new_n658), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n885), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n875), .A2(new_n752), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(KEYINPUT59), .A3(new_n883), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n884), .B1(new_n901), .B2(new_n903), .ZN(G1345gat));
  OAI21_X1  g703(.A(G155gat), .B1(new_n875), .B2(new_n888), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n882), .A2(new_n707), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n888), .A2(G155gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(G1346gat));
  NOR2_X1   g707(.A1(new_n848), .A2(new_n212), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n882), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n212), .B1(new_n875), .B2(new_n568), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n830), .A2(new_n665), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n832), .A2(new_n668), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT123), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n728), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n734), .A2(KEYINPUT124), .A3(new_n455), .A4(new_n668), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n732), .A2(new_n668), .A3(new_n733), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n773), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n919), .A2(new_n443), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n829), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n630), .A2(new_n293), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n917), .B2(new_n658), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n752), .B1(new_n324), .B2(new_n326), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n924), .B2(new_n928), .ZN(G1349gat));
  NAND3_X1  g728(.A1(new_n917), .A2(new_n304), .A3(new_n599), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n924), .A2(new_n599), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G183gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n923), .A2(new_n685), .A3(new_n829), .ZN(new_n938));
  INV_X1    g737(.A(G190gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n938), .B(new_n940), .C1(KEYINPUT125), .C2(KEYINPUT61), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n913), .A2(new_n303), .A3(new_n685), .A4(new_n915), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT126), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n886), .A2(new_n892), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n921), .A2(new_n676), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n950), .A2(new_n951), .A3(new_n630), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n676), .A2(new_n443), .A3(new_n707), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n913), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n728), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n952), .A2(new_n956), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n752), .A2(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n913), .A2(new_n953), .A3(new_n958), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  NAND3_X1  g759(.A1(new_n948), .A2(new_n658), .A3(new_n949), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n220), .A3(new_n599), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n599), .A3(new_n949), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n221), .A3(new_n685), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n949), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n971), .A2(new_n685), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n973), .B2(new_n221), .ZN(G1355gat));
endmodule


