//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n217), .ZN(new_n253));
  INV_X1    g0053(.A(G107), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n254), .A2(KEYINPUT23), .A3(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT23), .B1(new_n254), .B2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G116), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n255), .A2(new_n256), .B1(G20), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n209), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT22), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT22), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n263), .A2(new_n264), .A3(new_n209), .A4(G87), .ZN(new_n265));
  AOI211_X1 g0065(.A(KEYINPUT24), .B(new_n258), .C1(new_n262), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT24), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(new_n258), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n253), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n208), .A2(G33), .ZN(new_n273));
  AND4_X1   g0073(.A1(new_n217), .A2(new_n272), .A3(new_n252), .A4(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n254), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT25), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(new_n272), .B2(G107), .ZN(new_n278));
  AOI22_X1  g0078(.A1(G107), .A2(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  OAI211_X1 g0085(.A(G250), .B(new_n285), .C1(new_n259), .C2(new_n260), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G294), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT81), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n283), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT81), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n208), .A2(G45), .ZN(new_n293));
  OR2_X1    g0093(.A1(KEYINPUT5), .A2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(KEYINPUT5), .A2(G41), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n281), .B2(new_n282), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT5), .B(G41), .ZN(new_n300));
  INV_X1    g0100(.A(new_n293), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n300), .A2(new_n301), .B1(new_n281), .B2(new_n282), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G264), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n292), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n290), .A2(new_n291), .B1(G264), .B2(new_n302), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n299), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n280), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(new_n311), .A3(new_n299), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n280), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT82), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n312), .ZN(new_n317));
  INV_X1    g0117(.A(new_n280), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT82), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n280), .A2(new_n306), .A3(new_n309), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT8), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G58), .ZN(new_n325));
  INV_X1    g0125(.A(G58), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(KEYINPUT8), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT69), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n209), .A2(G33), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(KEYINPUT8), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(G58), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G20), .A2(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G150), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(KEYINPUT70), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n203), .A2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT70), .B1(new_n335), .B2(new_n337), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n253), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n253), .C1(new_n340), .C2(new_n341), .ZN(new_n345));
  INV_X1    g0145(.A(G50), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n275), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n252), .B(new_n217), .C1(G1), .C2(new_n209), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n343), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n298), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n283), .A2(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(G226), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n263), .A2(G222), .A3(new_n285), .ZN(new_n358));
  INV_X1    g0158(.A(G77), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n263), .A2(G1698), .ZN(new_n360));
  INV_X1    g0160(.A(G223), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n358), .B1(new_n359), .B2(new_n263), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(G169), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n308), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n351), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n351), .A2(KEYINPUT9), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT9), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n343), .A2(new_n370), .A3(new_n345), .A4(new_n350), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n364), .A2(new_n313), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G190), .B2(new_n364), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n374), .ZN(new_n376));
  AOI211_X1 g0176(.A(KEYINPUT10), .B(new_n376), .C1(new_n369), .C2(new_n371), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n367), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n253), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n330), .A2(G77), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n336), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT11), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n383), .A2(KEYINPUT11), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n385), .A2(KEYINPUT74), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT74), .B1(new_n385), .B2(new_n386), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT12), .B1(new_n272), .B2(G68), .ZN(new_n390));
  INV_X1    g0190(.A(new_n348), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n389), .A2(new_n390), .B1(new_n391), .B2(G68), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(G238), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n355), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n397), .A2(new_n399), .B1(new_n298), .B2(new_n353), .ZN(new_n400));
  OAI211_X1 g0200(.A(G232), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(new_n285), .C1(new_n259), .C2(new_n260), .ZN(new_n402));
  INV_X1    g0202(.A(G33), .ZN(new_n403));
  INV_X1    g0203(.A(G97), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n401), .B(new_n402), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n363), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n395), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(G238), .A3(new_n396), .ZN(new_n408));
  AND4_X1   g0208(.A1(new_n395), .A2(new_n406), .A3(new_n354), .A4(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n394), .B(G169), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n354), .A3(new_n408), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n400), .A2(new_n395), .A3(new_n406), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(G179), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n413), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n394), .B1(new_n416), .B2(G169), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n393), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n393), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(G200), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n311), .C2(new_n416), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n334), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n272), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n328), .A2(new_n334), .A3(new_n348), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n259), .A2(new_n260), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n428), .B2(new_n209), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT3), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n403), .ZN(new_n431));
  NAND2_X1  g0231(.A1(KEYINPUT3), .A2(G33), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n326), .A2(new_n221), .ZN(new_n436));
  OAI21_X1  g0236(.A(G20), .B1(new_n436), .B2(new_n202), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n336), .A2(G159), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT16), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n431), .A2(new_n209), .A3(new_n432), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT7), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n221), .B1(new_n444), .B2(new_n433), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n437), .A2(KEYINPUT16), .A3(new_n438), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n253), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n427), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G223), .B(new_n285), .C1(new_n259), .C2(new_n260), .ZN(new_n449));
  OAI211_X1 g0249(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G87), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n363), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n283), .A2(G232), .A3(new_n352), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n354), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n455), .A3(G179), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n354), .A2(new_n454), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n363), .B2(new_n452), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n305), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n448), .A2(KEYINPUT18), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n448), .A2(KEYINPUT75), .A3(KEYINPUT18), .A4(new_n459), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT18), .ZN(new_n464));
  INV_X1    g0264(.A(new_n459), .ZN(new_n465));
  INV_X1    g0265(.A(new_n427), .ZN(new_n466));
  INV_X1    g0266(.A(new_n446), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n380), .B1(new_n435), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT16), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n445), .B2(new_n439), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n466), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n464), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n462), .A2(new_n463), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n453), .A2(new_n455), .A3(G190), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n458), .B2(new_n313), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT17), .B1(new_n476), .B2(new_n471), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT17), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n448), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n275), .A2(new_n359), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n359), .B2(new_n348), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n331), .A2(new_n332), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n336), .B1(G20), .B2(G77), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT15), .B(G87), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n329), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n487), .B2(new_n253), .ZN(new_n488));
  INV_X1    g0288(.A(G244), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n354), .B1(new_n355), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n263), .A2(G232), .A3(new_n285), .ZN(new_n491));
  OAI221_X1 g0291(.A(new_n491), .B1(new_n254), .B2(new_n263), .C1(new_n360), .C2(new_n222), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n363), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n488), .B1(new_n493), .B2(new_n313), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n494), .A2(KEYINPUT72), .B1(G190), .B2(new_n493), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n488), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n493), .B2(G169), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n493), .A2(new_n308), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n422), .A2(new_n481), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n379), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT80), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(new_n285), .C1(new_n259), .C2(new_n260), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n431), .A2(G303), .A3(new_n432), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n511), .A2(new_n363), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n300), .A2(new_n301), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G270), .A3(new_n283), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n299), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT78), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n302), .A2(G270), .B1(new_n298), .B2(new_n296), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n363), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT78), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n209), .C1(G33), .C2(new_n404), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G20), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n253), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n522), .A2(KEYINPUT20), .A3(new_n253), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n272), .B2(G116), .ZN(new_n531));
  INV_X1    g0331(.A(G13), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(G1), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(KEYINPUT79), .A3(G20), .A4(new_n523), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n274), .A2(G116), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n305), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n516), .A2(new_n520), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n529), .A2(new_n535), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n517), .A2(new_n518), .A3(G179), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n516), .A2(KEYINPUT21), .A3(new_n520), .A4(new_n536), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n517), .A2(new_n519), .A3(new_n518), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n519), .B1(new_n517), .B2(new_n518), .ZN(new_n546));
  OAI21_X1  g0346(.A(G190), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n516), .A2(G200), .A3(new_n520), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n547), .A2(new_n540), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n507), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n543), .A2(new_n542), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n540), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT80), .A4(new_n539), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n263), .A2(G238), .A3(new_n285), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(new_n257), .C1(new_n360), .C2(new_n489), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n363), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n363), .A2(new_n301), .A3(new_n224), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n298), .B2(new_n301), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n305), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n263), .A2(new_n209), .A3(G68), .ZN(new_n562));
  NAND3_X1  g0362(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n209), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n206), .B2(G87), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n329), .A2(new_n404), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n562), .B(new_n565), .C1(KEYINPUT19), .C2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n253), .B1(new_n275), .B2(new_n486), .ZN(new_n568));
  INV_X1    g0368(.A(new_n274), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(new_n486), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n561), .B(new_n570), .C1(G179), .C2(new_n560), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n274), .A2(G87), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n560), .A2(G200), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n557), .A2(G190), .A3(new_n559), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n404), .A2(new_n254), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n205), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n254), .A2(KEYINPUT6), .A3(G97), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(G20), .B1(G77), .B2(new_n336), .ZN(new_n583));
  OAI21_X1  g0383(.A(G107), .B1(new_n429), .B2(new_n434), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n380), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n275), .A2(new_n404), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n569), .C2(new_n404), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G244), .B(new_n285), .C1(new_n259), .C2(new_n260), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT4), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(KEYINPUT77), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n593), .A2(new_n521), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n363), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n302), .A2(G257), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n299), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n590), .B1(new_n305), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n597), .B2(new_n363), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n308), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(G190), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n590), .C1(new_n313), .C2(new_n604), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n577), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n323), .A2(new_n506), .A3(new_n554), .A4(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n472), .A2(new_n460), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n421), .A2(new_n501), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n418), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n468), .A2(new_n470), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n453), .A2(new_n455), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n614), .A2(new_n427), .A3(new_n474), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n478), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n476), .A2(KEYINPUT17), .A3(new_n471), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n611), .B1(new_n613), .B2(new_n620), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n621), .A2(KEYINPUT84), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n375), .A2(new_n377), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n621), .B2(KEYINPUT84), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n622), .A2(new_n624), .B1(new_n351), .B2(new_n366), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n321), .B(KEYINPUT83), .ZN(new_n626));
  INV_X1    g0426(.A(new_n544), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n319), .A2(new_n577), .A3(new_n606), .A4(new_n608), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n571), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n577), .A2(KEYINPUT26), .A3(new_n605), .A4(new_n603), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n571), .A2(new_n576), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n606), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n625), .B1(new_n505), .B2(new_n638), .ZN(G369));
  NAND2_X1  g0439(.A1(new_n533), .A2(new_n209), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G213), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n554), .B1(new_n540), .B2(new_n646), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n627), .A2(new_n540), .A3(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G330), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n280), .A2(new_n645), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n323), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT85), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n323), .A2(KEYINPUT85), .A3(new_n654), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n321), .A2(new_n646), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n627), .A2(new_n645), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n657), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n626), .A2(new_n645), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n662), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n212), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n215), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  AOI211_X1 g0474(.A(KEYINPUT29), .B(new_n645), .C1(new_n630), .C2(new_n636), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n310), .A2(new_n544), .A3(KEYINPUT87), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT87), .B1(new_n310), .B2(new_n544), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n629), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(KEYINPUT86), .B2(new_n636), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n646), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n675), .B1(new_n681), .B2(KEYINPUT29), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n323), .A2(new_n554), .A3(new_n609), .A4(new_n646), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n560), .A2(new_n541), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n307), .A3(new_n604), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n684), .A2(KEYINPUT30), .A3(new_n604), .A4(new_n307), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n545), .A2(new_n546), .ZN(new_n689));
  AOI21_X1  g0489(.A(G179), .B1(new_n557), .B2(new_n559), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n602), .A3(new_n304), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n645), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT31), .B1(new_n692), .B2(new_n645), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n683), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n682), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n674), .B1(new_n699), .B2(G1), .ZN(G364));
  NAND2_X1  g0500(.A1(new_n650), .A2(new_n651), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n532), .A2(G20), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n208), .B1(new_n702), .B2(G45), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n669), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n701), .A2(new_n653), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n217), .B1(G20), .B2(new_n305), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n209), .A2(new_n308), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n311), .A3(new_n313), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n209), .A2(G190), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(G179), .A3(G200), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(G77), .A2(new_n712), .B1(new_n715), .B2(G68), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n313), .B2(G179), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n308), .A2(KEYINPUT90), .A3(G200), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n713), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G159), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT89), .B(KEYINPUT32), .Z(new_n725));
  OAI221_X1 g0525(.A(new_n716), .B1(new_n254), .B2(new_n720), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n718), .A2(new_n719), .A3(G20), .A4(G190), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n428), .B1(new_n728), .B2(G87), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(KEYINPUT91), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n724), .A2(new_n725), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n710), .A2(G190), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n313), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G50), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n732), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G58), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n209), .B1(new_n721), .B2(G190), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G97), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n731), .A2(new_n734), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n726), .A2(new_n730), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(KEYINPUT91), .B2(new_n729), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n733), .A2(G326), .ZN(new_n743));
  INV_X1    g0543(.A(new_n735), .ZN(new_n744));
  INV_X1    g0544(.A(G322), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(G294), .B2(new_n738), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT33), .B(G317), .Z(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n714), .B1(new_n711), .B2(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n263), .B(new_n750), .C1(G329), .C2(new_n723), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n727), .B(KEYINPUT92), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G303), .ZN(new_n753));
  INV_X1    g0553(.A(new_n720), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G283), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n747), .A2(new_n751), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n709), .B1(new_n742), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n708), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n668), .A2(new_n428), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G355), .B1(new_n523), .B2(new_n668), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n212), .A2(new_n428), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT88), .Z(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n215), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n250), .A2(G45), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n706), .B(new_n757), .C1(new_n761), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n760), .B(KEYINPUT93), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n649), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n707), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  AOI21_X1  g0573(.A(new_n645), .B1(new_n630), .B2(new_n636), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n501), .A2(new_n646), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n495), .A2(new_n496), .B1(new_n498), .B2(new_n645), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(new_n776), .B2(new_n501), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n774), .B(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n651), .B1(new_n683), .B2(new_n695), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n706), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(new_n782), .B2(KEYINPUT96), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(KEYINPUT96), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n708), .A2(new_n758), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n706), .B1(new_n359), .B2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G159), .A2(new_n712), .B1(new_n715), .B2(G150), .ZN(new_n787));
  INV_X1    g0587(.A(G137), .ZN(new_n788));
  INV_X1    g0588(.A(new_n733), .ZN(new_n789));
  INV_X1    g0589(.A(G143), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n787), .B1(new_n788), .B2(new_n789), .C1(new_n790), .C2(new_n744), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT34), .ZN(new_n792));
  INV_X1    g0592(.A(new_n752), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n791), .A2(new_n792), .B1(new_n346), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n720), .A2(new_n221), .ZN(new_n796));
  INV_X1    g0596(.A(G132), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n263), .B1(new_n737), .B2(new_n326), .C1(new_n797), .C2(new_n722), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n739), .B1(new_n749), .B2(new_n722), .C1(new_n744), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n711), .A2(new_n523), .B1(new_n714), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G303), .B2(new_n733), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT94), .Z(new_n805));
  AOI211_X1 g0605(.A(new_n801), .B(new_n805), .C1(G87), .C2(new_n754), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n263), .B1(new_n752), .B2(G107), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n775), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n497), .B1(new_n488), .B2(new_n646), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n502), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n786), .B1(new_n809), .B2(new_n709), .C1(new_n812), .C2(new_n759), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n784), .A2(new_n813), .ZN(G384));
  OR2_X1    g0614(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n815), .A2(G116), .A3(new_n218), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT36), .Z(new_n818));
  OAI211_X1 g0618(.A(new_n216), .B(G77), .C1(new_n326), .C2(new_n221), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n201), .A2(G68), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n208), .B(G13), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n418), .A2(new_n645), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT101), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT102), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT98), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n472), .A2(new_n463), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n620), .B1(new_n828), .B2(new_n462), .ZN(new_n829));
  INV_X1    g0629(.A(new_n643), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT97), .B1(new_n435), .B2(new_n440), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(KEYINPUT16), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n435), .A2(KEYINPUT97), .A3(new_n440), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n447), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n834), .B2(new_n466), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n827), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n481), .A2(KEYINPUT98), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT100), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n615), .A2(G169), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n614), .A2(new_n427), .B1(new_n842), .B2(new_n456), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT99), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n448), .A2(new_n844), .A3(new_n459), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n448), .A2(new_n830), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n617), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n840), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n448), .A2(new_n459), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT37), .B1(new_n850), .B2(KEYINPUT99), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n448), .A2(new_n475), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n643), .B1(new_n614), .B2(new_n427), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n851), .A2(new_n854), .A3(KEYINPUT100), .A4(new_n846), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n834), .A2(new_n466), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n459), .A2(new_n830), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n617), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n839), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT98), .B1(new_n481), .B2(new_n837), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n827), .B(new_n835), .C1(new_n473), .C2(new_n480), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n861), .B(KEYINPUT38), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT39), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n841), .B1(new_n854), .B2(new_n850), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n849), .B2(new_n855), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n847), .B1(new_n480), .B2(new_n611), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n865), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n826), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n869), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n868), .B1(new_n877), .B2(new_n865), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n865), .A2(new_n868), .A3(new_n873), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT102), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n825), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n611), .A2(new_n830), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n811), .A2(new_n502), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n810), .B1(new_n774), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n393), .A2(new_n645), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n418), .A2(new_n421), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n418), .B2(new_n421), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n877), .A2(new_n865), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n881), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n625), .B1(new_n682), .B2(new_n505), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n812), .B1(new_n886), .B2(new_n887), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n683), .B2(new_n695), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n862), .B2(new_n866), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n865), .A2(new_n873), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n900), .A3(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n506), .A2(new_n696), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(G330), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n208), .B2(new_n702), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n894), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n822), .B1(new_n908), .B2(new_n909), .ZN(G367));
  AND2_X1   g0710(.A1(new_n606), .A2(new_n608), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n645), .B1(new_n585), .B2(new_n589), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n603), .A2(new_n605), .A3(new_n645), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n657), .A2(new_n658), .A3(new_n663), .A4(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n911), .A2(new_n310), .A3(new_n912), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n645), .B1(new_n918), .B2(new_n606), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n916), .B2(KEYINPUT42), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI211_X1 g0722(.A(KEYINPUT103), .B(new_n919), .C1(new_n916), .C2(KEYINPUT42), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT104), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n573), .A2(new_n646), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n631), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n634), .B2(new_n926), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT43), .Z(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n917), .B(new_n931), .C1(new_n922), .C2(new_n923), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n924), .B2(new_n929), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT105), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n929), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT104), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT105), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(new_n938), .A3(new_n932), .A4(new_n930), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n662), .ZN(new_n941));
  INV_X1    g0741(.A(new_n915), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n666), .B2(new_n942), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n915), .B(new_n948), .C1(new_n664), .C2(new_n665), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n666), .B2(new_n942), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n664), .A2(KEYINPUT45), .A3(new_n665), .A4(new_n915), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n941), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n941), .B1(new_n950), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n661), .B1(new_n627), .B2(new_n645), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n959), .A2(new_n653), .A3(new_n664), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n653), .B1(new_n959), .B2(new_n664), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n698), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n669), .B(KEYINPUT41), .Z(new_n964));
  OAI21_X1  g0764(.A(new_n703), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n935), .A2(new_n943), .A3(new_n939), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n945), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n237), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n765), .ZN(new_n969));
  INV_X1    g0769(.A(new_n761), .ZN(new_n970));
  INV_X1    g0770(.A(new_n486), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n668), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n706), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n737), .A2(new_n221), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n789), .A2(new_n790), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(G150), .C2(new_n735), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n728), .A2(G58), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n754), .A2(G77), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n711), .A2(new_n201), .B1(new_n722), .B2(new_n788), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n428), .B(new_n979), .C1(G159), .C2(new_n715), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n789), .A2(new_n749), .B1(new_n737), .B2(new_n254), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G303), .B2(new_n735), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n752), .A2(KEYINPUT46), .A3(G116), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n727), .B2(new_n523), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n428), .B1(new_n711), .B2(new_n802), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n714), .A2(new_n800), .B1(new_n722), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n720), .A2(new_n404), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n983), .A2(new_n984), .A3(new_n986), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n981), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  OAI221_X1 g0794(.A(new_n973), .B1(new_n770), .B2(new_n928), .C1(new_n994), .C2(new_n709), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n967), .A2(new_n995), .ZN(G387));
  NAND2_X1  g0796(.A1(new_n962), .A2(new_n704), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n659), .A2(new_n660), .A3(new_n770), .ZN(new_n998));
  INV_X1    g0798(.A(new_n671), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n762), .A2(new_n999), .B1(new_n254), .B2(new_n668), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n484), .A2(new_n346), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT50), .Z(new_n1002));
  AOI21_X1  g0802(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n671), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n765), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G45), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n241), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1000), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n706), .B1(new_n1008), .B2(new_n761), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n263), .B1(new_n723), .B2(G326), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n727), .A2(new_n800), .B1(new_n802), .B2(new_n737), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G303), .A2(new_n712), .B1(new_n715), .B2(G311), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n988), .B2(new_n744), .C1(new_n745), .C2(new_n789), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1010), .B1(new_n523), .B2(new_n720), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n328), .A2(new_n334), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1020), .A2(new_n714), .B1(new_n221), .B2(new_n711), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT108), .ZN(new_n1022));
  INV_X1    g0822(.A(G150), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n263), .B1(new_n722), .B2(new_n1023), .C1(new_n744), .C2(new_n346), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n738), .A2(new_n971), .ZN(new_n1025));
  INV_X1    g0825(.A(G159), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n789), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n727), .A2(new_n359), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1024), .A2(new_n1027), .A3(new_n990), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1019), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1009), .B1(new_n1030), .B2(new_n709), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n962), .A2(new_n699), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n699), .B1(new_n960), .B2(new_n961), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n669), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n997), .B1(new_n998), .B2(new_n1031), .C1(new_n1032), .C2(new_n1034), .ZN(G393));
  NAND2_X1  g0835(.A1(new_n950), .A2(new_n954), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n662), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT109), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n955), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n956), .A2(KEYINPUT109), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1033), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT111), .A4(new_n1033), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1033), .A2(new_n957), .A3(new_n956), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n670), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n704), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n942), .A2(new_n760), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT110), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n247), .A2(new_n765), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n970), .B1(G97), .B2(new_n668), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n706), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n727), .A2(new_n802), .B1(new_n720), .B2(new_n254), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n715), .A2(G303), .B1(new_n723), .B2(G322), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n428), .C1(new_n800), .C2(new_n711), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(G116), .C2(new_n738), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n735), .A2(G311), .B1(new_n733), .B2(G317), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n712), .A2(new_n484), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n201), .B2(new_n714), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n737), .A2(new_n359), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n263), .B1(new_n722), .B2(new_n790), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n727), .A2(new_n221), .B1(new_n720), .B2(new_n223), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n735), .A2(G159), .B1(new_n733), .B2(G150), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT51), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n1059), .A2(new_n1061), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1052), .B(new_n1055), .C1(new_n709), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1050), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1048), .A2(new_n1073), .ZN(G390));
  NAND2_X1  g0874(.A1(new_n506), .A2(new_n779), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n625), .B(new_n1075), .C1(new_n682), .C2(new_n505), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT112), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n812), .B1(new_n697), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n888), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n697), .A2(new_n777), .A3(new_n888), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n646), .B(new_n883), .C1(new_n679), .C2(new_n680), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1083), .A2(new_n775), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n884), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n886), .B(new_n887), .C1(new_n779), .C2(new_n812), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n1081), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1076), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n867), .A2(new_n826), .A3(new_n874), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT102), .B1(new_n878), .B2(new_n879), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n824), .B1(new_n884), .B2(new_n888), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n824), .B(new_n900), .C1(new_n1084), .C2(new_n888), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n1082), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1082), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1090), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1081), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1094), .A2(new_n1095), .A3(new_n1082), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n1101), .A3(new_n1089), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(new_n669), .A3(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1091), .A2(new_n1092), .A3(new_n758), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n744), .A2(new_n797), .B1(new_n737), .B2(new_n1026), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G128), .B2(new_n733), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n714), .A2(new_n788), .B1(new_n722), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n428), .B(new_n1109), .C1(new_n712), .C2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1107), .B(new_n1112), .C1(new_n201), .C2(new_n720), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n728), .A2(G150), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT53), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n789), .A2(new_n802), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1064), .B(new_n1117), .C1(G116), .C2(new_n735), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n711), .A2(new_n404), .B1(new_n714), .B2(new_n254), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n428), .B1(new_n722), .B2(new_n800), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1119), .A2(new_n796), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1121), .C1(new_n223), .C2(new_n793), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n709), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n706), .B(new_n1123), .C1(new_n1020), .C2(new_n785), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1104), .A2(new_n704), .B1(new_n1105), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1103), .A2(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(KEYINPUT120), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n885), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n422), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n418), .A2(new_n421), .A3(new_n885), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n777), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n696), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n877), .B2(new_n865), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n901), .C1(new_n1133), .C2(KEYINPUT40), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n351), .A2(new_n830), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT118), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n378), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n367), .B(new_n1137), .C1(new_n375), .C2(new_n377), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1139), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT119), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1134), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT119), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1139), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1148), .A2(new_n899), .A3(G330), .A4(new_n901), .ZN(new_n1149));
  AND4_X1   g0949(.A1(new_n881), .A2(new_n1145), .A3(new_n891), .A4(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n881), .A2(new_n891), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1127), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n892), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n881), .A2(new_n1145), .A3(new_n891), .A4(new_n1149), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT120), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1076), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1102), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1076), .B1(new_n1104), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT57), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n669), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n758), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(G33), .A2(G41), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT113), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT116), .B(G124), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n722), .A2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G159), .C2(new_n754), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n733), .A2(G125), .B1(G150), .B2(new_n738), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n744), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n711), .A2(new_n788), .B1(new_n714), .B2(new_n797), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT115), .Z(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(new_n728), .C2(new_n1111), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1172), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1179), .B2(new_n1178), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n789), .A2(new_n523), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n974), .B(new_n1182), .C1(G107), .C2(new_n735), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n720), .A2(new_n326), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT114), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n711), .A2(new_n486), .B1(new_n714), .B2(new_n404), .ZN(new_n1186));
  INV_X1    g0986(.A(G41), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(new_n428), .C1(new_n722), .C2(new_n802), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1186), .A2(new_n1028), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT58), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1169), .B(new_n346), .C1(G41), .C2(new_n263), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n708), .B1(new_n1181), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n706), .B1(new_n201), .B2(new_n785), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT117), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1167), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1157), .B2(new_n704), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1166), .A2(new_n1201), .ZN(G375));
  INV_X1    g1002(.A(new_n964), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1085), .A2(new_n1076), .A3(new_n1088), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1090), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n888), .A2(new_n758), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1025), .B1(new_n789), .B2(new_n800), .C1(new_n802), .C2(new_n744), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n712), .A2(G107), .B1(new_n723), .B2(G303), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n263), .B1(new_n715), .B2(G116), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1209), .A2(new_n978), .A3(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(new_n404), .C2(new_n793), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n263), .B1(new_n722), .B2(new_n1174), .C1(new_n711), .C2(new_n1023), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G50), .B2(new_n738), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n1185), .C1(new_n1026), .C2(new_n793), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT121), .Z(new_n1216));
  AOI22_X1  g1016(.A1(new_n733), .A2(G132), .B1(new_n715), .B2(new_n1111), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n788), .B2(new_n744), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1212), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1219), .A2(new_n708), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n706), .B(new_n1220), .C1(new_n221), .C2(new_n785), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1161), .A2(new_n704), .B1(new_n1206), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1205), .A2(new_n1222), .ZN(G381));
  NOR4_X1   g1023(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1072), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1225));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OR3_X1    g1027(.A1(G375), .A2(new_n1227), .A3(G387), .ZN(G407));
  INV_X1    g1028(.A(G375), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n644), .A3(new_n1226), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(new_n1230), .A3(G213), .ZN(G409));
  XNOR2_X1  g1031(.A(G393), .B(new_n772), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT123), .B1(G387), .B2(new_n1225), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G387), .A2(new_n1225), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G387), .A2(KEYINPUT123), .A3(new_n1225), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT125), .B1(G387), .B2(new_n1225), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(G390), .A2(new_n1239), .A3(new_n995), .A4(new_n967), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G387), .A2(KEYINPUT124), .A3(new_n1225), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT124), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1232), .B1(new_n1234), .B2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1232), .A2(new_n1237), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(G343), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1201), .C1(new_n1160), .C2(new_n1165), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1150), .A2(new_n1151), .A3(new_n1127), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT120), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1159), .B(new_n1203), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1200), .B1(new_n1163), .B2(new_n704), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1226), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1247), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1204), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1090), .B2(KEYINPUT60), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1085), .A2(new_n1076), .A3(new_n1088), .A4(KEYINPUT60), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n669), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1222), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n784), .A3(new_n813), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G384), .B(new_n1222), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1247), .A2(G2897), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1264), .B(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1247), .B(new_n1264), .C1(new_n1248), .C2(new_n1254), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1247), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1264), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1245), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1271), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1265), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1264), .B(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1278), .B(new_n1279), .C1(new_n1255), .C2(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(KEYINPUT122), .B(KEYINPUT63), .C1(new_n1255), .C2(new_n1273), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT122), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1274), .B2(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1282), .A2(new_n1283), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1237), .A2(new_n1232), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1277), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(KEYINPUT122), .B1(new_n1269), .B2(KEYINPUT63), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1274), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1292), .A2(new_n1267), .A3(new_n1293), .A4(new_n1278), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1294), .A2(new_n1245), .A3(KEYINPUT126), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1276), .B1(new_n1291), .B2(new_n1295), .ZN(G405));
  NOR2_X1   g1096(.A1(new_n1229), .A2(G378), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1248), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1264), .A2(KEYINPUT127), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1264), .A2(KEYINPUT127), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1245), .A2(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1288), .A2(new_n1289), .A3(new_n1302), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1301), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1290), .A2(KEYINPUT127), .A3(new_n1264), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1245), .A2(new_n1302), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1300), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(G402));
endmodule


