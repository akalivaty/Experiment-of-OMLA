//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT68), .A2(G119), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT68), .A2(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n195), .B2(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(G128), .B1(new_n193), .B2(new_n194), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n196), .B1(new_n201), .B2(new_n192), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT76), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n212), .A2(KEYINPUT76), .A3(G140), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n211), .B2(KEYINPUT16), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT77), .A4(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n208), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT79), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n223), .B(new_n208), .C1(new_n216), .C2(new_n220), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n218), .A2(new_n219), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n212), .A2(KEYINPUT76), .A3(G140), .ZN(new_n227));
  XNOR2_X1  g041(.A(G125), .B(G140), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(KEYINPUT76), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(G146), .C1(new_n209), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n216), .A2(new_n220), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT78), .A3(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n207), .B1(new_n225), .B2(new_n235), .ZN(new_n236));
  OR3_X1    g050(.A1(new_n201), .A2(KEYINPUT80), .A3(new_n205), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT80), .B1(new_n201), .B2(new_n205), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n237), .B(new_n238), .C1(new_n202), .C2(G110), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n208), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n239), .A2(new_n230), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n191), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT78), .B1(new_n233), .B2(G146), .ZN(new_n244));
  NOR4_X1   g058(.A1(new_n216), .A2(new_n220), .A3(new_n231), .A4(new_n208), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n222), .B(new_n224), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n207), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n230), .A3(new_n240), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n190), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n242), .A2(new_n250), .A3(KEYINPUT25), .A4(new_n243), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G217), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(G234), .B2(new_n243), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n255), .A2(KEYINPUT81), .A3(new_n257), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n242), .A2(new_n250), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n257), .A2(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n198), .B2(G116), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n195), .B2(G116), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n198), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT68), .A2(G119), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n271), .A2(KEYINPUT69), .A3(G116), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n266), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n276));
  INV_X1    g090(.A(G113), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT67), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(KEYINPUT2), .B2(G113), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n278), .A2(new_n280), .B1(KEYINPUT2), .B2(G113), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n271), .A2(G116), .A3(new_n272), .ZN(new_n283));
  INV_X1    g097(.A(new_n268), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n273), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n275), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n273), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n281), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n208), .A2(G143), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G146), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT0), .A4(G128), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G143), .B(G146), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n297), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT0), .B(G128), .Z(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT11), .B1(new_n305), .B2(G137), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G137), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G134), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n306), .A2(new_n309), .B1(new_n305), .B2(G137), .ZN(new_n310));
  INV_X1    g124(.A(G131), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n299), .A2(new_n313), .A3(new_n302), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n304), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  AOI21_X1  g130(.A(G128), .B1(new_n291), .B2(new_n293), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n292), .A2(KEYINPUT1), .A3(G146), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(KEYINPUT66), .B(new_n318), .C1(new_n297), .C2(G128), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n297), .A2(new_n322), .A3(G128), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n310), .A2(new_n311), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n308), .B2(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n305), .B2(G137), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n326), .A2(new_n308), .A3(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(G131), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n290), .A2(new_n315), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n287), .A2(new_n289), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n299), .A2(new_n313), .A3(new_n302), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n313), .B1(new_n299), .B2(new_n302), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n310), .B(G131), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n331), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n333), .B1(new_n341), .B2(new_n332), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n332), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n290), .B1(new_n331), .B2(new_n315), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n188), .A3(G210), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT27), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G101), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n344), .A2(new_n348), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n315), .A2(KEYINPUT30), .A3(new_n331), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n331), .B1(new_n338), .B2(new_n303), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n335), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n332), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n354), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(KEYINPUT74), .A3(new_n354), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n332), .A2(new_n333), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n359), .A2(new_n335), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n290), .A2(new_n315), .A3(KEYINPUT28), .A4(new_n331), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n355), .B1(new_n372), .B2(new_n354), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n243), .B(new_n357), .C1(new_n368), .C2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n362), .A2(new_n353), .A3(new_n332), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT31), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n362), .A2(KEYINPUT31), .A3(new_n353), .A4(new_n332), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n377), .A2(new_n378), .B1(new_n354), .B2(new_n372), .ZN(new_n379));
  NOR2_X1   g193(.A1(G472), .A2(G902), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT72), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n374), .A2(G472), .B1(KEYINPUT32), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n377), .A2(new_n378), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n372), .A2(new_n354), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n387));
  INV_X1    g201(.A(new_n381), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT73), .B1(new_n379), .B2(new_n381), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT32), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n265), .B1(new_n383), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G214), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G104), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(G107), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n397), .A2(G107), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n400), .A2(G104), .ZN(new_n406));
  OAI21_X1  g220(.A(G101), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n289), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G113), .B1(new_n283), .B2(KEYINPUT5), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n288), .B2(KEYINPUT5), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n275), .B2(new_n286), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n289), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n404), .A2(new_n407), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n418), .B(KEYINPUT8), .Z(new_n419));
  OAI21_X1  g233(.A(KEYINPUT87), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n273), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT70), .B1(new_n285), .B2(new_n273), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT5), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n410), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n409), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G101), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n427), .B(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n425), .A2(new_n426), .B1(new_n335), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT86), .B1(new_n324), .B2(G125), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n303), .A2(G125), .ZN(new_n433));
  AND4_X1   g247(.A1(new_n322), .A2(new_n291), .A3(new_n293), .A4(G128), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n318), .B1(new_n297), .B2(G128), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n316), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n212), .A4(new_n321), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT7), .B1(new_n440), .B2(G953), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n431), .A2(new_n418), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n420), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n444));
  INV_X1    g258(.A(new_n419), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n408), .B1(new_n425), .B2(new_n289), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n444), .B(new_n445), .C1(new_n446), .C2(new_n412), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n433), .A2(new_n438), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n449));
  INV_X1    g263(.A(new_n441), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n432), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT88), .B1(new_n439), .B2(new_n441), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(KEYINPUT89), .B(new_n243), .C1(new_n443), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n431), .B2(new_n418), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n418), .B2(new_n431), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n440), .A2(G953), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n439), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n431), .ZN(new_n461));
  INV_X1    g275(.A(new_n418), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n420), .A2(new_n442), .A3(new_n447), .A4(new_n453), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT89), .B1(new_n466), .B2(new_n243), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n396), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT91), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n243), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(KEYINPUT90), .A3(new_n464), .A4(new_n455), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n470), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n476), .A3(new_n464), .A4(new_n455), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n395), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT9), .B(G234), .Z(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT82), .ZN(new_n480));
  OAI21_X1  g294(.A(G221), .B1(new_n480), .B2(G902), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT83), .Z(new_n482));
  INV_X1    g296(.A(G469), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n243), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n408), .B1(new_n435), .B2(new_n434), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n320), .A2(new_n416), .A3(new_n321), .A4(new_n323), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n486), .A2(KEYINPUT85), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n436), .A2(new_n489), .A3(new_n321), .A4(new_n416), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n312), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n486), .A2(KEYINPUT85), .A3(new_n487), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n493), .A2(KEYINPUT12), .A3(new_n312), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n430), .A2(new_n304), .A3(new_n314), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT10), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n416), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n486), .A2(new_n497), .B1(new_n324), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n499), .A3(new_n338), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G110), .B(G140), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n188), .A2(G227), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT84), .Z(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n496), .A2(new_n499), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n312), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n501), .A2(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n484), .B1(new_n510), .B2(G469), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n500), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n504), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n495), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n483), .A3(new_n243), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n482), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G113), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n397), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT19), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n214), .B2(new_n215), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n228), .A2(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n208), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n230), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n522), .B1(new_n230), .B2(new_n526), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n349), .A2(new_n188), .A3(G214), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n292), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n349), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n311), .A3(new_n531), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n527), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT18), .A2(G131), .ZN(new_n537));
  OR3_X1    g351(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n532), .B2(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n229), .A2(G146), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n240), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n521), .B1(new_n536), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n532), .A2(KEYINPUT17), .A3(G131), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n520), .B(new_n543), .C1(new_n246), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(G475), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n557), .A3(new_n552), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n225), .A2(new_n235), .A3(new_n548), .A4(new_n547), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n520), .B1(new_n559), .B2(new_n543), .ZN(new_n560));
  INV_X1    g374(.A(new_n550), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n243), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n556), .A2(new_n558), .B1(G475), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n188), .A2(G952), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n480), .A2(new_n256), .A3(G953), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n575));
  INV_X1    g389(.A(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(KEYINPUT95), .A2(G122), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G116), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n576), .A2(G116), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G116), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n577), .B2(new_n578), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT96), .B1(new_n586), .B2(new_n582), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n584), .A2(new_n587), .A3(G107), .ZN(new_n588));
  AOI21_X1  g402(.A(G107), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n292), .A2(G128), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT13), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n292), .B2(G128), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n199), .A2(KEYINPUT97), .A3(G143), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(KEYINPUT98), .A3(G134), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n596), .A2(new_n591), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n305), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n305), .B1(new_n592), .B2(new_n596), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n590), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n589), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n583), .A2(KEYINPUT14), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n583), .A2(KEYINPUT14), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n580), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G107), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n600), .A2(new_n305), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n596), .A2(new_n591), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G134), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n605), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n574), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n609), .A3(new_n613), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(new_n573), .C1(new_n590), .C2(new_n603), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G478), .ZN(new_n619));
  NOR2_X1   g433(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  AOI211_X1 g439(.A(G902), .B(new_n623), .C1(new_n615), .C2(new_n617), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n563), .A2(KEYINPUT100), .A3(new_n572), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n552), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n545), .B2(new_n550), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n558), .B1(new_n554), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n562), .A2(G475), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n627), .A3(new_n572), .A4(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n518), .B1(new_n628), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n393), .A2(new_n478), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT101), .B(G101), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G3));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n394), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n477), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n465), .A2(new_n467), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n395), .B1(new_n643), .B2(new_n476), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n470), .B1(new_n465), .B2(new_n467), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n640), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n615), .A2(new_n617), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT33), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n615), .A2(new_n650), .A3(new_n617), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(G478), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n618), .A2(new_n619), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n619), .A2(new_n243), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n563), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n647), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n260), .A2(new_n517), .A3(new_n261), .A4(new_n264), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n379), .B2(G902), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n389), .A2(new_n390), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n572), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NAND2_X1  g480(.A1(new_n630), .A2(new_n554), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n556), .A2(new_n667), .B1(G475), .B2(new_n562), .ZN(new_n668));
  INV_X1    g482(.A(new_n627), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n644), .A2(new_n646), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n643), .A2(new_n640), .A3(new_n394), .A4(new_n476), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n572), .A3(new_n663), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NAND2_X1  g490(.A1(new_n248), .A2(new_n249), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n677), .B(new_n678), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n263), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n260), .A2(new_n261), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n662), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n478), .A3(new_n636), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  NAND2_X1  g499(.A1(new_n382), .A2(KEYINPUT32), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n357), .A2(new_n243), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT74), .B1(new_n363), .B2(new_n354), .ZN(new_n688));
  AOI211_X1 g502(.A(new_n365), .B(new_n353), .C1(new_n362), .C2(new_n332), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n373), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n392), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n511), .A2(new_n516), .ZN(new_n693));
  INV_X1    g507(.A(new_n482), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n568), .A2(G900), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n566), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT81), .B1(new_n255), .B2(new_n257), .ZN(new_n698));
  INV_X1    g512(.A(new_n257), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n259), .B(new_n699), .C1(new_n253), .C2(new_n254), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n697), .B1(new_n701), .B2(new_n680), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n692), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n673), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  NAND2_X1  g519(.A1(new_n475), .A2(new_n477), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT38), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n260), .A2(new_n261), .A3(new_n680), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n709), .A2(new_n395), .A3(new_n563), .A4(new_n627), .ZN(new_n710));
  INV_X1    g524(.A(G472), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n345), .A2(new_n346), .A3(new_n353), .ZN(new_n712));
  AOI211_X1 g526(.A(G902), .B(new_n712), .C1(new_n353), .C2(new_n363), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n392), .B(new_n686), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n696), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n517), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n710), .A2(new_n714), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n708), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n292), .ZN(G45));
  NAND2_X1  g535(.A1(new_n659), .A2(new_n703), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NAND2_X1  g537(.A1(new_n515), .A2(new_n243), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n516), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n482), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n393), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n473), .A2(new_n464), .A3(new_n455), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT102), .B1(new_n729), .B2(new_n470), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n477), .A2(new_n394), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n672), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n572), .A3(new_n657), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT41), .B(G113), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  INV_X1    g550(.A(new_n670), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n572), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n728), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT103), .B(G116), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G18));
  AOI22_X1  g555(.A1(new_n635), .A2(new_n628), .B1(new_n701), .B2(new_n680), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n732), .A3(new_n692), .A4(new_n727), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  OAI211_X1 g558(.A(new_n343), .B(KEYINPUT28), .C1(new_n345), .C2(new_n346), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n369), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n342), .A2(new_n343), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n354), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n384), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n388), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n661), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n265), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n563), .A2(new_n627), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n726), .A2(new_n482), .A3(new_n571), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n732), .A2(new_n752), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  NAND2_X1  g570(.A1(new_n386), .A2(new_n243), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n757), .A2(G472), .B1(new_n749), .B2(new_n388), .ZN(new_n758));
  INV_X1    g572(.A(new_n696), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n563), .A2(new_n656), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n709), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n732), .A3(new_n727), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT104), .ZN(new_n764));
  INV_X1    g578(.A(new_n727), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n671), .B2(new_n672), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n762), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n475), .A2(new_n394), .A3(new_n477), .A4(new_n517), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n391), .B1(new_n379), .B2(new_n381), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n691), .A2(new_n686), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n264), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n698), .A2(new_n700), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n777), .A3(new_n760), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n771), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n692), .A2(new_n777), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n760), .A2(new_n771), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n772), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT105), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n475), .A2(new_n394), .A3(new_n477), .ZN(new_n784));
  INV_X1    g598(.A(new_n781), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n393), .A3(new_n517), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n775), .A2(new_n777), .A3(new_n760), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT42), .B1(new_n787), .B2(new_n772), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT105), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n311), .ZN(G33));
  NOR2_X1   g606(.A1(new_n670), .A2(new_n759), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n784), .A2(new_n393), .A3(new_n517), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT106), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n773), .A2(new_n796), .A3(new_n393), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n510), .A2(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n509), .A2(new_n506), .A3(new_n500), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n496), .A2(new_n499), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n804), .A2(new_n338), .B1(new_n492), .B2(new_n494), .ZN(new_n805));
  INV_X1    g619(.A(new_n505), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n483), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT107), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n802), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g625(.A(KEYINPUT107), .B(new_n483), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT108), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(G469), .B1(new_n510), .B2(KEYINPUT45), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT107), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n810), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n802), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n801), .B(new_n484), .C1(new_n813), .C2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(G469), .B(G902), .C1(new_n513), .C2(new_n514), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n800), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n813), .A2(new_n818), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n801), .B1(new_n823), .B2(new_n484), .ZN(new_n824));
  INV_X1    g638(.A(new_n484), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(KEYINPUT46), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(KEYINPUT109), .A3(new_n516), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n694), .A3(new_n715), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n630), .A2(new_n554), .ZN(new_n831));
  AOI211_X1 g645(.A(KEYINPUT20), .B(new_n629), .C1(new_n545), .C2(new_n550), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n632), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n656), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n631), .A2(KEYINPUT110), .A3(new_n632), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n833), .A2(new_n656), .A3(KEYINPUT43), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n662), .A3(new_n709), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT44), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n475), .A2(new_n394), .A3(new_n477), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n840), .B1(new_n838), .B2(KEYINPUT43), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT44), .A3(new_n662), .A4(new_n709), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n844), .A2(new_n845), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT112), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n846), .B(KEYINPUT111), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n844), .A4(new_n850), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n830), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G137), .ZN(G39));
  NAND2_X1  g672(.A1(new_n265), .A2(new_n760), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n846), .A2(new_n692), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n828), .A2(KEYINPUT47), .A3(new_n694), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT47), .B1(new_n828), .B2(new_n694), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(G140), .ZN(G42));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n846), .A2(new_n765), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n714), .A2(new_n265), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n567), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n868), .A2(new_n833), .A3(new_n836), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n849), .A2(new_n567), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n866), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n681), .A3(new_n751), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n708), .A2(new_n395), .A3(new_n727), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n708), .A2(new_n876), .A3(new_n395), .A4(new_n727), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n870), .A2(new_n752), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n861), .A2(new_n862), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n694), .B2(new_n726), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n853), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT115), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n865), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n880), .B(new_n881), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n888), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT51), .A4(new_n873), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n265), .B(new_n871), .C1(new_n383), .C2(new_n774), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n879), .A2(new_n766), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n564), .C1(new_n658), .C2(new_n868), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n890), .A2(new_n893), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n703), .B(new_n732), .C1(new_n657), .C2(new_n737), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n709), .A2(new_n697), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n732), .A2(new_n714), .A3(new_n902), .A4(new_n753), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n767), .B1(new_n766), .B2(new_n762), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n647), .A2(new_n761), .A3(KEYINPUT104), .A4(new_n765), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n901), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT52), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n769), .A2(KEYINPUT52), .A3(new_n901), .A4(new_n903), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n789), .B1(new_n786), .B2(new_n788), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n728), .B1(new_n733), .B2(new_n738), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n563), .A2(new_n627), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n915), .B(new_n572), .C1(new_n563), .C2(new_n836), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n478), .A2(new_n663), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n743), .A2(new_n755), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n637), .A2(new_n683), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n772), .A2(new_n761), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT113), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n668), .A2(new_n627), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n703), .A2(new_n923), .A3(new_n784), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n692), .A2(new_n702), .A3(new_n925), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT113), .B1(new_n927), .B2(new_n846), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n922), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n913), .A2(new_n921), .A3(new_n798), .A4(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT53), .B1(new_n910), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n798), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n743), .A2(new_n755), .A3(new_n918), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n637), .A2(new_n683), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n692), .A2(new_n777), .A3(new_n727), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n572), .B(new_n935), .C1(new_n659), .C2(new_n673), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n932), .A2(new_n791), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT114), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT53), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT114), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n906), .A2(new_n941), .A3(new_n907), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n931), .A2(new_n943), .A3(KEYINPUT54), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n940), .B1(new_n910), .B2(new_n930), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT54), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n786), .A2(new_n788), .A3(KEYINPUT53), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n932), .A2(new_n937), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n939), .A3(new_n942), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n900), .A2(new_n951), .B1(G952), .B2(G953), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n395), .B(new_n482), .C1(new_n726), .C2(KEYINPUT49), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(KEYINPUT49), .B2(new_n726), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n838), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n708), .A2(new_n867), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(G75));
  NAND2_X1  g771(.A1(new_n945), .A2(new_n949), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(G902), .A3(new_n470), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT56), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n458), .A2(new_n463), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n460), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT55), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n959), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n959), .B2(new_n960), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n188), .A2(G952), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(G51));
  NAND3_X1  g782(.A1(new_n958), .A2(G902), .A3(new_n823), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT119), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n484), .B(KEYINPUT57), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n946), .B1(new_n945), .B2(new_n949), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n515), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n967), .B1(new_n970), .B2(new_n975), .ZN(G54));
  AND2_X1   g790(.A1(KEYINPUT58), .A2(G475), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n948), .A2(new_n939), .A3(new_n942), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n908), .A2(new_n909), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT53), .B1(new_n938), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(G902), .B(new_n977), .C1(new_n978), .C2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n545), .A3(new_n550), .ZN(new_n982));
  INV_X1    g796(.A(new_n967), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n958), .A2(G902), .A3(new_n551), .A4(new_n977), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT120), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT120), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n982), .A2(new_n987), .A3(new_n983), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G60));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n649), .A2(new_n651), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT121), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n654), .B(KEYINPUT59), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT54), .B1(new_n978), .B2(new_n980), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n950), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n990), .B1(new_n997), .B2(new_n967), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n994), .B1(new_n972), .B2(new_n973), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(KEYINPUT122), .A3(new_n983), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n944), .A2(new_n950), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n992), .B1(new_n1001), .B2(new_n993), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n998), .A2(new_n1000), .A3(new_n1002), .ZN(G63));
  NAND2_X1  g817(.A1(G217), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT60), .Z(new_n1005));
  NAND2_X1  g819(.A1(new_n958), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n262), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n958), .A2(new_n679), .A3(new_n1005), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1008), .A2(new_n983), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT61), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n983), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(G66));
  OAI21_X1  g828(.A(G953), .B1(new_n570), .B2(new_n440), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n921), .B2(G953), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n961), .B1(G898), .B2(new_n188), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT123), .Z(new_n1018));
  XNOR2_X1  g832(.A(new_n1016), .B(new_n1018), .ZN(G69));
  NAND2_X1  g833(.A1(new_n769), .A2(new_n901), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1020), .B1(new_n830), .B2(new_n856), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n732), .A2(new_n777), .A3(new_n753), .A4(new_n775), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n829), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1021), .A2(new_n863), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n798), .A2(new_n783), .A3(new_n790), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT125), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT125), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n913), .A2(new_n1028), .A3(new_n798), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(KEYINPUT126), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n829), .B1(new_n852), .B2(new_n855), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n1032), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT126), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1033), .A2(new_n1034), .A3(new_n863), .A4(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1031), .A2(new_n1036), .A3(new_n188), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n358), .A2(new_n361), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n524), .A2(new_n525), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  AOI21_X1  g854(.A(new_n1040), .B1(G900), .B2(G953), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT124), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n769), .B(new_n901), .C1(new_n708), .C2(new_n719), .ZN(new_n1044));
  OR2_X1    g858(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n915), .B1(new_n563), .B2(new_n836), .ZN(new_n1046));
  NOR4_X1   g860(.A1(new_n780), .A2(new_n846), .A3(new_n716), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1047), .B1(new_n1044), .B2(KEYINPUT62), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n1045), .A2(new_n1048), .A3(new_n857), .A4(new_n863), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n188), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1043), .B1(new_n1050), .B2(new_n1040), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1042), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1053), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1042), .A2(new_n1055), .A3(new_n1051), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1054), .A2(new_n1056), .ZN(G72));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  OAI21_X1  g873(.A(new_n1059), .B1(new_n1049), .B2(new_n937), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1060), .A2(new_n353), .A3(new_n363), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n931), .A2(new_n943), .ZN(new_n1062));
  INV_X1    g876(.A(new_n375), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n1063), .B1(new_n368), .B2(KEYINPUT127), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1064), .B1(KEYINPUT127), .B2(new_n368), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1065), .A2(new_n1059), .ZN(new_n1066));
  OAI211_X1 g880(.A(new_n1061), .B(new_n983), .C1(new_n1062), .C2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n1031), .A2(new_n1036), .A3(new_n921), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1068), .A2(new_n1059), .ZN(new_n1069));
  NOR2_X1   g883(.A1(new_n363), .A2(new_n353), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(G57));
endmodule


