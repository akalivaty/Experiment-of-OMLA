//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT70), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(new_n190), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(G104), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n203), .A2(G107), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n203), .A2(G107), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n201), .A2(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n197), .A3(KEYINPUT69), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(KEYINPUT2), .B2(G113), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n214), .A2(new_n216), .B1(KEYINPUT2), .B2(G113), .ZN(new_n217));
  INV_X1    g031(.A(new_n191), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n199), .A2(new_n212), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G101), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n224), .A3(G101), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n217), .B1(new_n192), .B2(new_n194), .ZN(new_n227));
  INV_X1    g041(.A(new_n219), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n220), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G110), .B(G122), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n220), .B(new_n231), .C1(new_n226), .C2(new_n229), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT6), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT0), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n236), .A2(KEYINPUT65), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT0), .A4(G128), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT77), .A2(G125), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT77), .A2(G125), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(KEYINPUT0), .B2(G128), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT64), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n239), .A2(new_n246), .A3(new_n249), .A4(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n254), .A2(KEYINPUT87), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT68), .B(G128), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(G143), .B2(new_n240), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n244), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n241), .A2(new_n243), .A3(new_n257), .A4(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n261), .A2(new_n249), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(KEYINPUT87), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G224), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n266), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n255), .A2(new_n263), .A3(new_n268), .A4(new_n262), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n230), .A2(new_n271), .A3(new_n232), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n235), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n254), .B(KEYINPUT87), .Z(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n268), .A4(new_n262), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT7), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n264), .B1(new_n277), .B2(new_n266), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n197), .B(new_n196), .C1(new_n218), .C2(KEYINPUT5), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n212), .B1(new_n279), .B2(new_n228), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n199), .A2(new_n211), .A3(new_n219), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n231), .B(KEYINPUT8), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n276), .A2(new_n278), .A3(new_n234), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n273), .A2(new_n274), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT88), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n273), .A2(new_n284), .A3(new_n274), .A4(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n211), .A2(new_n259), .A3(new_n260), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT84), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n236), .A2(new_n296), .A3(new_n257), .A4(G128), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n244), .B1(new_n258), .B2(new_n238), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n294), .B1(new_n299), .B2(new_n211), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT11), .ZN(new_n302));
  INV_X1    g116(.A(G137), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .A4(G134), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n305), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n303), .B2(G134), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G131), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n306), .B2(new_n304), .ZN(new_n314));
  INV_X1    g128(.A(G131), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(G131), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND4_X1   g132(.A1(KEYINPUT12), .A2(new_n300), .A3(new_n313), .A4(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n318), .A2(new_n313), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT12), .B1(new_n320), .B2(new_n300), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT85), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n212), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n318), .A2(new_n313), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n239), .A2(new_n246), .A3(new_n253), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n223), .A2(new_n328), .A3(new_n225), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n212), .A2(KEYINPUT10), .A3(new_n261), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n327), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G140), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G227), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n337));
  INV_X1    g151(.A(new_n300), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(new_n327), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n300), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n322), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n320), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n331), .ZN(new_n346));
  INV_X1    g160(.A(new_n335), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G469), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n274), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n274), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n331), .B1(new_n319), .B2(new_n321), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n353), .A2(new_n347), .B1(new_n336), .B2(new_n345), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n354), .B2(G469), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT9), .B(G234), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G221), .B1(new_n358), .B2(G902), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n359), .B(KEYINPUT81), .Z(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT82), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n293), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  AOI211_X1 g177(.A(KEYINPUT86), .B(new_n361), .C1(new_n351), .C2(new_n355), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n291), .B(new_n292), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G237), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n333), .A3(G214), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT89), .B(G143), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n371), .B2(new_n242), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G131), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT18), .ZN(new_n376));
  OAI21_X1  g190(.A(G140), .B1(new_n247), .B2(new_n248), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G140), .C1(new_n247), .C2(new_n248), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT76), .B1(new_n381), .B2(G140), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n383));
  INV_X1    g197(.A(G140), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G125), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G146), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(G140), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n240), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT18), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n370), .B(new_n372), .C1(new_n393), .C2(new_n315), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT90), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(KEYINPUT90), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n376), .A2(new_n392), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(KEYINPUT19), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT19), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(KEYINPUT19), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n400), .A2(new_n389), .A3(new_n390), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n240), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n386), .A4(new_n380), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n249), .A2(new_n405), .A3(new_n384), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(G146), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(KEYINPUT92), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n370), .A2(new_n315), .A3(new_n372), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n374), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT92), .B1(new_n403), .B2(new_n407), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n397), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G113), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n203), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n375), .A2(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n404), .A2(new_n406), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n240), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT17), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n374), .A2(new_n421), .A3(new_n409), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n418), .A2(new_n420), .A3(new_n407), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n397), .A3(new_n415), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(KEYINPUT93), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n427));
  INV_X1    g241(.A(new_n402), .ZN(new_n428));
  AOI211_X1 g242(.A(G146), .B(new_n428), .C1(new_n387), .C2(KEYINPUT19), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n404), .A2(G146), .A3(new_n406), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n408), .A3(new_n410), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n415), .B1(new_n432), .B2(new_n397), .ZN(new_n433));
  INV_X1    g247(.A(new_n424), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n426), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT20), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n433), .B2(new_n434), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G475), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n415), .B1(new_n423), .B2(new_n397), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n444), .B2(new_n274), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n438), .A2(new_n441), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n333), .A2(G952), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(G234), .B2(G237), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT96), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT21), .B(G898), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n449), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  INV_X1    g273(.A(G122), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G116), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT94), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n201), .B1(new_n462), .B2(KEYINPUT14), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(G116), .B2(new_n460), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n463), .B(new_n464), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n256), .A2(G143), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n238), .B2(G143), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT95), .B(G134), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n305), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(new_n467), .Z(new_n473));
  XNOR2_X1  g287(.A(new_n464), .B(G107), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n357), .A2(G217), .A3(new_n333), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n459), .B1(new_n482), .B2(G902), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n481), .B(new_n274), .C1(KEYINPUT15), .C2(new_n458), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n447), .A2(new_n457), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT97), .B1(new_n365), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n292), .ZN(new_n489));
  AOI211_X1 g303(.A(G469), .B(G902), .C1(new_n343), .C2(new_n348), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n353), .A2(new_n347), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n336), .A2(new_n345), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(G469), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n352), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n362), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT86), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n356), .A2(new_n293), .A3(new_n362), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n489), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n438), .A2(new_n441), .A3(new_n446), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n500), .A2(new_n456), .A3(new_n485), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT97), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(new_n291), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n488), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n256), .A2(G119), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(G119), .B2(new_n238), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT24), .B(G110), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT75), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n187), .B2(G128), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n512), .C1(G119), .C2(new_n238), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n508), .B1(new_n513), .B2(G110), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n391), .A3(new_n407), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(G110), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n420), .A2(new_n407), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n516), .B(new_n517), .C1(new_n506), .C2(new_n507), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT22), .B(G137), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n518), .A3(new_n522), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n274), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n527));
  INV_X1    g341(.A(G217), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(G234), .B2(new_n274), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n524), .A2(new_n530), .A3(new_n274), .A4(new_n525), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n529), .A2(G902), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n525), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT79), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n534), .A2(KEYINPUT79), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n318), .A2(new_n328), .A3(new_n313), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n303), .A2(G134), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n305), .A2(G137), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n261), .B(new_n543), .C1(G131), .C2(new_n311), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n540), .A2(new_n229), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT30), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n548), .A3(new_n544), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n229), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT31), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT26), .B(G101), .Z(new_n554));
  NAND3_X1  g368(.A1(new_n366), .A2(new_n333), .A3(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n556), .B(new_n557), .Z(new_n558));
  NAND4_X1  g372(.A1(new_n552), .A2(KEYINPUT72), .A3(new_n553), .A4(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n540), .A2(new_n548), .A3(new_n544), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n548), .B1(new_n540), .B2(new_n544), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n551), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n540), .A2(new_n229), .A3(new_n544), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n562), .A2(KEYINPUT72), .A3(new_n563), .A4(new_n558), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n229), .B1(new_n540), .B2(new_n544), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT28), .B1(new_n545), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT28), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n558), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n559), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(G472), .A2(G902), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n573), .A2(KEYINPUT32), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT32), .B1(new_n573), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n229), .B1(new_n547), .B2(new_n549), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n571), .B1(new_n578), .B2(new_n545), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT29), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n567), .A2(new_n569), .A3(new_n558), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT73), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n581), .A2(new_n580), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G902), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n579), .A2(new_n586), .A3(new_n580), .A4(new_n581), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n539), .B1(new_n577), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n573), .A2(new_n574), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT32), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n573), .A2(KEYINPUT32), .A3(new_n574), .ZN(new_n594));
  AND4_X1   g408(.A1(new_n539), .A2(new_n589), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n538), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT80), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT74), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n577), .A2(new_n539), .A3(new_n589), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n537), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n504), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT98), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G3));
  NOR2_X1   g420(.A1(new_n363), .A2(new_n364), .ZN(new_n607));
  INV_X1    g421(.A(new_n286), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n285), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n290), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n292), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT99), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n613), .A3(new_n292), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n457), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n591), .ZN(new_n616));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n573), .B2(new_n274), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NOR4_X1   g433(.A1(new_n607), .A2(new_n615), .A3(new_n619), .A4(new_n537), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n621));
  OR2_X1    g435(.A1(new_n481), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n481), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n622), .A2(G478), .A3(new_n624), .A4(new_n274), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n458), .B1(new_n482), .B2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n500), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n437), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n425), .B2(new_n435), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n445), .B1(new_n634), .B2(KEYINPUT20), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT93), .B1(new_n417), .B2(new_n424), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n433), .A2(new_n426), .A3(new_n434), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n437), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n440), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n620), .A2(new_n485), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  INV_X1    g457(.A(new_n619), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n519), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n533), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n532), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n504), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  INV_X1    g465(.A(new_n449), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(new_n452), .B2(G900), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n635), .A2(new_n639), .A3(new_n485), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n600), .A2(new_n601), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n612), .A2(new_n614), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n648), .B1(new_n363), .B2(new_n364), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n656), .A2(new_n657), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XOR2_X1   g477(.A(new_n653), .B(KEYINPUT39), .Z(new_n664));
  NOR2_X1   g478(.A1(new_n607), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n447), .B(new_n486), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n578), .A2(new_n545), .A3(new_n571), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n545), .A2(new_n566), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n668), .B1(new_n670), .B2(new_n571), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n577), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n665), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n674), .B1(new_n675), .B2(KEYINPUT40), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n291), .A2(KEYINPUT38), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n291), .A2(KEYINPUT38), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n648), .A2(new_n489), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n667), .A2(new_n676), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND3_X1  g497(.A1(new_n500), .A2(new_n627), .A3(new_n653), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n657), .A2(new_n659), .A3(new_n661), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND2_X1  g501(.A1(new_n349), .A2(new_n274), .ZN(new_n688));
  AND2_X1   g502(.A1(KEYINPUT102), .A2(G469), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n360), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n615), .A2(new_n628), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n657), .A2(new_n694), .A3(new_n538), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NOR3_X1   g511(.A1(new_n537), .A2(new_n693), .A3(new_n456), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(new_n485), .A3(new_n640), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n658), .B1(new_n600), .B2(new_n601), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  INV_X1    g520(.A(new_n648), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n487), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n693), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n657), .A2(new_n708), .A3(new_n659), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NOR3_X1   g525(.A1(new_n658), .A2(new_n447), .A3(new_n486), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n574), .A2(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n574), .A2(KEYINPUT104), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n573), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n618), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n712), .A2(new_n698), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AND2_X1   g532(.A1(new_n716), .A2(new_n648), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n658), .A2(new_n693), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n685), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  OAI21_X1  g536(.A(new_n691), .B1(new_n490), .B2(new_n495), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n291), .A2(new_n489), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n356), .A2(new_n726), .A3(new_n691), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n684), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(new_n538), .C1(new_n590), .C2(new_n595), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n599), .A2(KEYINPUT42), .A3(new_n538), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n730), .A2(new_n731), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n315), .ZN(G33));
  INV_X1    g548(.A(new_n728), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n602), .A2(new_n656), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n619), .A2(new_n648), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT107), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT43), .B1(new_n447), .B2(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n447), .A2(new_n627), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n447), .B(new_n627), .C1(KEYINPUT106), .C2(KEYINPUT43), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n739), .A2(KEYINPUT44), .A3(new_n744), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n725), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n354), .A2(KEYINPUT45), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n354), .A2(KEYINPUT45), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(G469), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n494), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n351), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT46), .B1(new_n754), .B2(new_n494), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n691), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(new_n664), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n747), .A2(KEYINPUT108), .A3(new_n725), .A4(new_n748), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n751), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  XNOR2_X1  g577(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n758), .B1(new_n766), .B2(KEYINPUT47), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n684), .A2(new_n538), .ZN(new_n769));
  INV_X1    g583(.A(new_n725), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n657), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n384), .ZN(G42));
  XOR2_X1   g587(.A(new_n628), .B(KEYINPUT111), .Z(new_n774));
  INV_X1    g588(.A(new_n365), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n619), .A2(new_n537), .A3(new_n456), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n604), .A2(KEYINPUT112), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n604), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n500), .A2(new_n486), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n649), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n778), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n730), .A2(new_n731), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n732), .A2(new_n729), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n729), .A2(new_n719), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n497), .A2(new_n498), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n788), .A2(new_n640), .A3(new_n648), .A4(new_n725), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n486), .A2(new_n653), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n657), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n736), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n723), .B1(new_n577), .B2(new_n672), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n712), .A2(new_n707), .A3(new_n653), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n662), .A2(new_n686), .A3(new_n721), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n721), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n658), .B(new_n660), .C1(new_n600), .C2(new_n601), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(new_n656), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT52), .A3(new_n686), .A4(new_n795), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n793), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n710), .A2(new_n695), .A3(new_n717), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n703), .B2(new_n704), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n597), .B(new_n537), .C1(new_n600), .C2(new_n601), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n488), .A2(new_n503), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n777), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n782), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n604), .A2(KEYINPUT112), .A3(new_n777), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n805), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n657), .A2(new_n656), .A3(new_n538), .A4(new_n735), .ZN(new_n818));
  INV_X1    g632(.A(new_n787), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n733), .A2(new_n818), .A3(new_n791), .A4(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n796), .A2(new_n797), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n796), .A2(new_n797), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n807), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n806), .A2(new_n824), .A3(KEYINPUT113), .ZN(new_n825));
  INV_X1    g639(.A(new_n817), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT53), .A4(new_n803), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n806), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n693), .A2(new_n770), .A3(new_n652), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n744), .A2(new_n599), .A3(new_n538), .A4(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT48), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n690), .A2(new_n692), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n362), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n765), .B2(new_n767), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n537), .A2(new_n652), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n744), .A2(new_n716), .A3(new_n725), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n652), .B(new_n537), .C1(new_n742), .C2(new_n743), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n679), .A2(KEYINPUT114), .A3(new_n489), .A4(new_n709), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n677), .A2(new_n489), .A3(new_n678), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n693), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n841), .A2(new_n846), .A3(KEYINPUT50), .A4(new_n716), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n744), .A2(new_n716), .A3(new_n838), .ZN(new_n849));
  INV_X1    g663(.A(new_n846), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n674), .A2(new_n838), .A3(new_n709), .A4(new_n725), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n447), .A3(new_n626), .A4(new_n625), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n744), .A2(new_n719), .A3(new_n832), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n855), .C1(new_n837), .C2(new_n839), .ZN(new_n856));
  OAI211_X1 g670(.A(KEYINPUT51), .B(new_n840), .C1(new_n852), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n856), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n840), .A2(KEYINPUT51), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n847), .A2(new_n851), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n448), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n841), .A2(new_n716), .A3(new_n720), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n853), .A2(new_n629), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n834), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n829), .A2(new_n831), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  OR2_X1    g681(.A1(G952), .A2(G953), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n829), .A2(new_n865), .A3(new_n869), .A4(new_n831), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n679), .B1(new_n873), .B2(KEYINPUT110), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n537), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n361), .B(new_n673), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n741), .B1(new_n873), .B2(KEYINPUT110), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n292), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(KEYINPUT117), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(G75));
  AND2_X1   g697(.A1(new_n235), .A2(new_n272), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(new_n270), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n806), .A2(new_n824), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n274), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n333), .A2(G952), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n886), .A2(new_n891), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n889), .B2(new_n288), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(G51));
  NAND2_X1  g710(.A1(new_n494), .A2(KEYINPUT57), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n494), .A2(KEYINPUT57), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n888), .A2(new_n830), .ZN(new_n899));
  INV_X1    g713(.A(new_n831), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n897), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n349), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n888), .A2(new_n274), .A3(new_n754), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n893), .B1(new_n902), .B2(new_n903), .ZN(G54));
  INV_X1    g718(.A(new_n893), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n906));
  INV_X1    g720(.A(new_n436), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT118), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n906), .A2(KEYINPUT118), .A3(new_n907), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G60));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n829), .B2(new_n831), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n622), .A2(new_n624), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n899), .B2(new_n900), .ZN(new_n920));
  OAI221_X1 g734(.A(new_n905), .B1(new_n918), .B2(new_n919), .C1(new_n920), .C2(new_n917), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(G63));
  XNOR2_X1  g736(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n528), .A2(new_n274), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n887), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n646), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n905), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n524), .A2(new_n525), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(new_n926), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g746(.A(G953), .B1(new_n455), .B2(new_n265), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n826), .B2(G953), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT121), .Z(new_n935));
  INV_X1    g749(.A(G898), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n884), .B1(new_n936), .B2(G953), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  NAND2_X1  g752(.A1(new_n398), .A2(new_n402), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT122), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n550), .B(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n760), .A2(new_n599), .A3(new_n538), .A4(new_n712), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n942), .A2(new_n786), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n762), .A2(new_n736), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n801), .A2(KEYINPUT123), .A3(new_n686), .ZN(new_n945));
  INV_X1    g759(.A(new_n772), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n662), .A2(new_n686), .A3(new_n721), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n952), .B2(new_n333), .ZN(new_n953));
  INV_X1    g767(.A(G900), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n954), .B2(G227), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n333), .B1(G227), .B2(G900), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n809), .A2(new_n810), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n774), .A2(new_n780), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n957), .A2(new_n665), .A3(new_n725), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n772), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n762), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n945), .A2(new_n682), .A3(new_n949), .ZN(new_n962));
  NOR2_X1   g776(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n956), .B1(new_n965), .B2(new_n333), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n953), .A2(new_n955), .B1(new_n966), .B2(new_n941), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n579), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n668), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT127), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n825), .A2(new_n828), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n552), .B(KEYINPUT125), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n961), .A2(new_n826), .A3(new_n964), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n969), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n558), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n976), .B2(new_n558), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n905), .B(new_n973), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n952), .A2(new_n826), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n558), .B1(new_n981), .B2(new_n969), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n974), .B2(new_n982), .ZN(G57));
endmodule


