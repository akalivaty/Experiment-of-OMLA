//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n191));
  OAI211_X1 g005(.A(G119), .B(new_n190), .C1(new_n191), .C2(KEYINPUT72), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n193), .B(KEYINPUT23), .C1(new_n194), .C2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G110), .ZN(new_n197));
  AOI22_X1  g011(.A1(KEYINPUT72), .A2(new_n191), .B1(new_n194), .B2(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G119), .B(G128), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(G146), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n202), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n201), .A2(new_n200), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n196), .A2(new_n198), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n204), .A2(G146), .A3(new_n207), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n204), .B2(new_n207), .ZN(new_n217));
  OAI221_X1 g031(.A(new_n214), .B1(new_n215), .B2(new_n197), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n202), .A2(KEYINPUT73), .A3(new_n208), .A4(new_n210), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XOR2_X1   g037(.A(new_n221), .B(new_n223), .Z(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n213), .A2(new_n218), .A3(new_n219), .A4(new_n224), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n188), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n189), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n226), .A2(new_n227), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n189), .A2(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT28), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT66), .B1(new_n242), .B2(G134), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n240), .A3(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n244), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n240), .A2(G137), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n242), .A2(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT64), .A2(G143), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT64), .A2(G143), .ZN(new_n255));
  OAI21_X1  g069(.A(G146), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n209), .A2(G143), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(new_n261), .A3(G128), .A4(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n258), .A3(new_n260), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT64), .A2(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n209), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n209), .A2(G143), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(G128), .A2(new_n265), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n250), .B(new_n253), .C1(new_n264), .C2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n254), .A2(new_n255), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n275), .B2(new_n209), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT0), .B(G128), .Z(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT65), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(new_n272), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n277), .ZN(new_n282));
  INV_X1    g096(.A(new_n262), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n268), .A2(new_n269), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G146), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT0), .A3(G128), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n246), .A2(new_n248), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n241), .A2(new_n243), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n288), .A2(G131), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n245), .B1(new_n244), .B2(new_n249), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n274), .B(KEYINPUT70), .C1(new_n287), .C2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT2), .B(G113), .Z(new_n294));
  XNOR2_X1  g108(.A(G116), .B(G119), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n294), .B(new_n295), .Z(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n250), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n279), .A3(new_n282), .A4(new_n286), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT70), .B1(new_n300), .B2(new_n274), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n238), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n274), .B(new_n296), .C1(new_n287), .C2(new_n292), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n300), .B2(new_n274), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n222), .A3(G210), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT69), .Z(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n274), .B1(new_n287), .B2(new_n292), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT30), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n296), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n300), .A2(KEYINPUT30), .A3(new_n274), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n303), .A2(new_n312), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n303), .A2(new_n323), .A3(new_n312), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT31), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT31), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n320), .A2(new_n322), .A3(new_n327), .A4(new_n324), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G472), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n188), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT71), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n329), .A2(new_n333), .A3(new_n330), .A4(new_n188), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT32), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n329), .A2(KEYINPUT32), .A3(new_n330), .A4(new_n188), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n302), .A2(new_n306), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n302), .A2(new_n306), .A3(new_n312), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n320), .A2(new_n303), .ZN(new_n341));
  INV_X1    g155(.A(new_n312), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n336), .B1(new_n344), .B2(new_n330), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n237), .B1(new_n335), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G475), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n308), .A2(new_n222), .A3(G143), .A4(G214), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n308), .A2(new_n222), .A3(G214), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT86), .B(new_n349), .C1(new_n275), .C2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n349), .A2(KEYINPUT86), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(new_n245), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT17), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n216), .A2(new_n217), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n308), .A2(new_n222), .A3(G214), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n284), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n352), .B1(new_n360), .B2(new_n349), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G131), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n245), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n356), .B(new_n357), .C1(new_n364), .C2(KEYINPUT17), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n203), .A2(new_n209), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n210), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n354), .A2(KEYINPUT87), .B1(KEYINPUT18), .B2(G131), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n369), .B(new_n370), .C1(new_n351), .C2(new_n353), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G113), .B(G122), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT90), .B(G104), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n376), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n365), .A2(new_n378), .A3(new_n372), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n348), .B1(new_n380), .B2(new_n188), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n367), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n370), .B1(new_n361), .B2(new_n369), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n354), .A2(KEYINPUT87), .A3(KEYINPUT18), .A4(G131), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT19), .B1(new_n203), .B2(KEYINPUT88), .ZN(new_n387));
  INV_X1    g201(.A(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G140), .ZN(new_n389));
  AND4_X1   g203(.A1(KEYINPUT88), .A2(new_n206), .A3(new_n389), .A4(KEYINPUT19), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n209), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n208), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n362), .B2(new_n363), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT89), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n391), .A2(new_n208), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n361), .A2(G131), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n355), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n372), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n399), .A3(new_n376), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n379), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT20), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n348), .A4(new_n188), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(G475), .B1(new_n400), .B2(new_n379), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n402), .B1(new_n405), .B2(new_n188), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n382), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT91), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n348), .A3(new_n188), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT20), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n382), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n267), .A2(G128), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n284), .B2(G128), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n416), .A2(new_n240), .ZN(new_n417));
  XNOR2_X1  g231(.A(G116), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G107), .ZN(new_n420));
  INV_X1    g234(.A(G107), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n284), .A2(G128), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(KEYINPUT13), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n423), .B1(new_n240), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G116), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT14), .A3(G122), .ZN(new_n429));
  OAI211_X1 g243(.A(G107), .B(new_n429), .C1(new_n419), .C2(KEYINPUT14), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n416), .A2(new_n240), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n422), .B(new_n430), .C1(new_n417), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT9), .B(G234), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n435), .A2(new_n187), .A3(G953), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n427), .A2(new_n432), .A3(new_n436), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT15), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n414), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G221), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n434), .B2(new_n188), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n188), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT74), .B1(new_n421), .B2(G104), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n453));
  INV_X1    g267(.A(G104), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(G107), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G101), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT3), .B1(new_n454), .B2(G107), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n421), .A3(G104), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n454), .A2(G107), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n421), .A2(G104), .ZN(new_n463));
  OAI21_X1  g277(.A(G101), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n190), .B1(new_n466), .B2(new_n262), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n263), .B1(new_n276), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT79), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n461), .A2(new_n464), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT77), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n190), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n263), .B1(new_n475), .B2(new_n285), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n465), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n465), .B2(new_n476), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n469), .B(new_n473), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n292), .A2(KEYINPUT78), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n479), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT81), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n477), .A2(new_n478), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n473), .A2(new_n469), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT12), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT10), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n470), .A2(new_n492), .A3(new_n472), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n458), .A2(new_n460), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n457), .B1(new_n494), .B2(new_n456), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n495), .A2(new_n496), .B1(new_n461), .B2(KEYINPUT4), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n452), .A2(new_n455), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n458), .A2(new_n460), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(G101), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT76), .B1(new_n503), .B2(new_n287), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n461), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n500), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n279), .A2(new_n282), .A3(new_n286), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT76), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n493), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n492), .B1(new_n477), .B2(new_n478), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n292), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G110), .B(G140), .ZN(new_n515));
  INV_X1    g329(.A(G227), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G953), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n515), .B(new_n517), .Z(new_n518));
  NAND4_X1  g332(.A1(new_n484), .A2(new_n491), .A3(new_n514), .A4(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n518), .ZN(new_n520));
  INV_X1    g334(.A(new_n493), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n510), .B1(new_n508), .B2(new_n509), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n513), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n299), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n299), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n519), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n451), .B1(new_n529), .B2(new_n450), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n488), .A2(new_n490), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n520), .B1(new_n531), .B2(new_n527), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n514), .A2(new_n525), .A3(new_n518), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n532), .A2(KEYINPUT80), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT80), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(G469), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n449), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n222), .A2(G952), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(G234), .B2(G237), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT21), .B(G898), .Z(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n188), .B(new_n222), .C1(G234), .C2(G237), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(G110), .B(G122), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n194), .A2(G116), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n428), .A2(G119), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT5), .ZN(new_n549));
  OR3_X1    g363(.A1(new_n428), .A2(KEYINPUT5), .A3(G119), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(G113), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n294), .A2(new_n295), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n472), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n546), .B(new_n555), .C1(new_n503), .C2(new_n296), .ZN(new_n556));
  INV_X1    g370(.A(new_n546), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n296), .B1(new_n506), .B2(new_n507), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n554), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n559), .A3(KEYINPUT6), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT6), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n561), .B(new_n557), .C1(new_n558), .C2(new_n554), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n287), .A2(G125), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n470), .A2(new_n388), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n287), .A2(KEYINPUT82), .A3(G125), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G224), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G953), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n566), .A2(new_n573), .A3(new_n567), .A4(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n563), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n546), .B(KEYINPUT8), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n461), .A2(new_n464), .B1(new_n551), .B2(new_n552), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n554), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT83), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT83), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(new_n580), .C1(new_n554), .C2(new_n581), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n564), .A2(new_n567), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n577), .B2(new_n571), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT84), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n579), .A2(new_n586), .A3(new_n588), .A4(KEYINPUT84), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n556), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G210), .B1(G237), .B2(G902), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n576), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n576), .B2(new_n593), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT85), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n576), .A2(new_n593), .A3(new_n594), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n543), .B(new_n545), .C1(new_n597), .C2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n347), .A2(new_n447), .A3(new_n537), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n332), .A2(new_n334), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n329), .A2(new_n188), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n530), .B2(new_n536), .ZN(new_n608));
  INV_X1    g422(.A(new_n543), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n576), .A2(new_n593), .ZN(new_n610));
  INV_X1    g424(.A(new_n594), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n545), .B1(new_n612), .B2(new_n598), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n236), .A2(new_n449), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n608), .A2(new_n609), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n438), .A2(new_n439), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(G478), .A3(new_n188), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n440), .A2(G478), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(KEYINPUT92), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(KEYINPUT92), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n414), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT34), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  INV_X1    g440(.A(new_n446), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n403), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n405), .A2(KEYINPUT93), .A3(new_n402), .A4(new_n188), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n410), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n382), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n615), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n220), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n234), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n232), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n607), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n641), .A2(new_n601), .A3(new_n447), .A4(new_n537), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(KEYINPUT32), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n604), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n345), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n613), .A2(new_n639), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n539), .B1(new_n542), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n632), .A2(new_n627), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n537), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT94), .ZN(new_n654));
  INV_X1    g468(.A(new_n449), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n519), .A2(new_n528), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n450), .A3(new_n188), .ZN(new_n657));
  INV_X1    g471(.A(new_n451), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT80), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n482), .A2(new_n483), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n518), .B1(new_n661), .B2(new_n514), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n514), .A2(new_n525), .A3(new_n518), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n532), .A2(KEYINPUT80), .A3(new_n533), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n450), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n655), .B1(new_n659), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n345), .B1(new_n604), .B2(new_n645), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT94), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n649), .A4(new_n652), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n654), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n414), .A2(new_n446), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n651), .B(KEYINPUT39), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n678), .B(new_n544), .C1(new_n677), .C2(new_n676), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n598), .A2(new_n599), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n612), .A2(new_n598), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(KEYINPUT85), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT38), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(new_n639), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n313), .B1(new_n304), .B2(new_n305), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n325), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n330), .B1(new_n686), .B2(new_n188), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n646), .A2(new_n336), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT95), .ZN(new_n690));
  INV_X1    g504(.A(new_n336), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n335), .A2(new_n691), .A3(new_n687), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n679), .A2(new_n684), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n284), .ZN(G45));
  INV_X1    g511(.A(new_n651), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n412), .B1(new_n411), .B2(new_n382), .ZN(new_n699));
  AOI211_X1 g513(.A(KEYINPUT91), .B(new_n381), .C1(new_n410), .C2(new_n403), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n622), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT96), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT96), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n414), .A2(new_n703), .A3(new_n622), .A4(new_n698), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n648), .A2(new_n537), .A3(new_n649), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n209), .ZN(G48));
  NAND2_X1  g522(.A1(new_n656), .A2(new_n188), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n655), .A2(new_n710), .A3(new_n613), .A4(new_n657), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n414), .A2(new_n609), .A3(new_n622), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n347), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NOR3_X1   g529(.A1(new_n632), .A2(new_n627), .A3(new_n543), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n711), .A2(new_n648), .A3(new_n237), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NOR2_X1   g532(.A1(new_n529), .A2(new_n450), .ZN(new_n719));
  AOI211_X1 g533(.A(G469), .B(G902), .C1(new_n519), .C2(new_n528), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n449), .A4(new_n543), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n648), .A2(new_n721), .A3(new_n447), .A4(new_n649), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AND3_X1   g537(.A1(new_n329), .A2(new_n330), .A3(new_n188), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n330), .B1(new_n329), .B2(new_n188), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n724), .A2(new_n725), .A3(new_n236), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n414), .A2(new_n726), .A3(new_n446), .A4(new_n613), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n721), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT97), .B(G122), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G24));
  NAND3_X1  g544(.A1(new_n606), .A2(new_n331), .A3(new_n639), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT98), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n606), .A2(KEYINPUT98), .A3(new_n331), .A4(new_n639), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n702), .A2(new_n711), .A3(new_n735), .A4(new_n704), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(new_n705), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n724), .A2(KEYINPUT32), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n237), .B1(new_n739), .B2(new_n345), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT99), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n662), .A2(new_n663), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n657), .A2(new_n743), .A3(new_n658), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n655), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n597), .A2(new_n544), .A3(new_n600), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n738), .A2(new_n741), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n346), .A2(new_n746), .A3(new_n745), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n748), .A2(KEYINPUT42), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  AND3_X1   g566(.A1(new_n347), .A2(new_n747), .A3(new_n652), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n240), .ZN(G36));
  INV_X1    g568(.A(KEYINPUT101), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n408), .A2(new_n622), .A3(new_n413), .ZN(new_n756));
  NAND2_X1  g570(.A1(KEYINPUT100), .A2(KEYINPUT43), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT100), .B(KEYINPUT43), .Z(new_n759));
  OAI21_X1  g573(.A(new_n758), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(new_n607), .A3(new_n639), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT44), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n597), .A2(new_n544), .A3(new_n600), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n755), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI211_X1 g578(.A(KEYINPUT101), .B(new_n746), .C1(new_n761), .C2(KEYINPUT44), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(KEYINPUT44), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n664), .A2(new_n768), .A3(new_n665), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(G469), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n658), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n658), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n657), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n655), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(new_n675), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT102), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n775), .A2(new_n657), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n771), .B2(new_n658), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n783), .B(new_n655), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n776), .B2(new_n655), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n787), .A2(new_n788), .A3(new_n705), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n668), .A3(new_n236), .A4(new_n763), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  INV_X1    g605(.A(KEYINPUT103), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n614), .A2(new_n544), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n683), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n719), .A2(new_n720), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT104), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n756), .B(new_n794), .C1(KEYINPUT49), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT105), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n792), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n799), .A3(new_n695), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n736), .B1(new_n706), .B2(new_n705), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n232), .A2(new_n638), .A3(new_n698), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT109), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n232), .A2(new_n808), .A3(new_n638), .A4(new_n698), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n744), .A2(new_n810), .A3(new_n655), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n414), .A2(new_n446), .A3(new_n613), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n689), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n811), .A2(new_n689), .A3(new_n812), .A4(KEYINPUT110), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n805), .A2(new_n672), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n805), .A2(new_n817), .A3(new_n672), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n713), .A2(new_n717), .A3(new_n722), .A4(new_n728), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT106), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n710), .A2(new_n613), .A3(new_n655), .A4(new_n657), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n346), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n826), .A2(new_n716), .B1(new_n721), .B2(new_n727), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT106), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n713), .A4(new_n722), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT107), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n446), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT107), .B1(new_n444), .B2(new_n445), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n413), .A3(new_n408), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n623), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n608), .A2(new_n836), .A3(new_n601), .A4(new_n614), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n747), .A2(new_n704), .A3(new_n702), .A4(new_n735), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n602), .A3(new_n838), .A4(new_n642), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n667), .A2(new_n668), .A3(new_n640), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n632), .A2(new_n651), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n832), .A2(new_n833), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n682), .A2(new_n544), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(KEYINPUT108), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n537), .B(new_n639), .C1(new_n335), .C2(new_n345), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n753), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n830), .A2(new_n751), .A3(new_n840), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n803), .B1(new_n822), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n749), .A2(new_n652), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT108), .B1(new_n841), .B2(new_n845), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n848), .A2(new_n847), .A3(new_n844), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT111), .B1(new_n857), .B2(new_n839), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(new_n850), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n823), .A2(new_n803), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n751), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n861), .A2(new_n821), .A3(new_n819), .A4(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n802), .A2(new_n852), .A3(new_n853), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n804), .B1(new_n671), .B2(new_n654), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n820), .B1(new_n866), .B2(new_n817), .ZN(new_n867));
  INV_X1    g681(.A(new_n821), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n857), .A2(new_n839), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(new_n751), .A3(new_n830), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n852), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n802), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n852), .A2(new_n853), .A3(new_n864), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n865), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n760), .A2(new_n539), .A3(new_n726), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n825), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n692), .B(KEYINPUT95), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n719), .A2(new_n720), .A3(new_n449), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n763), .A2(KEYINPUT116), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n710), .A2(new_n655), .A3(new_n657), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n746), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n885), .A3(new_n237), .A4(new_n539), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT118), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n882), .A2(new_n885), .A3(new_n539), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n695), .A4(new_n237), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n414), .A2(new_n622), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n760), .A2(new_n539), .A3(new_n882), .A4(new_n885), .ZN(new_n893));
  INV_X1    g707(.A(new_n735), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT117), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n888), .A2(new_n896), .A3(new_n735), .A4(new_n760), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT51), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n892), .A2(new_n900), .A3(new_n898), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT50), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n881), .A2(KEYINPUT113), .A3(new_n545), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n710), .A2(new_n655), .A3(new_n657), .A4(new_n545), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n683), .A2(new_n908), .A3(KEYINPUT114), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT114), .B1(new_n683), .B2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n878), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n903), .B1(new_n911), .B2(KEYINPUT115), .ZN(new_n912));
  INV_X1    g726(.A(new_n910), .ZN(new_n913));
  INV_X1    g727(.A(new_n878), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n683), .A2(new_n908), .A3(KEYINPUT114), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT50), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n787), .A2(new_n788), .B1(new_n655), .B2(new_n796), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n763), .A3(new_n914), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n902), .A2(new_n912), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT120), .B1(new_n901), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n912), .A2(new_n918), .A3(new_n920), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n892), .A2(new_n898), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(KEYINPUT119), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n923), .A2(new_n924), .A3(new_n927), .A4(new_n902), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n888), .A2(new_n741), .A3(new_n760), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT48), .ZN(new_n931));
  AND4_X1   g745(.A1(new_n414), .A2(new_n887), .A3(new_n890), .A4(new_n622), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n899), .A2(new_n918), .A3(new_n912), .A4(new_n920), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n538), .B(new_n932), .C1(new_n933), .C2(new_n925), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n877), .A2(new_n879), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(G952), .A2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n801), .B1(new_n936), .B2(new_n937), .ZN(G75));
  NOR2_X1   g752(.A1(new_n222), .A2(G952), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n188), .B1(new_n852), .B2(new_n864), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT56), .B1(new_n941), .B2(G210), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n560), .A2(new_n562), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n575), .B(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n948), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(G51));
  NAND2_X1  g765(.A1(new_n658), .A2(KEYINPUT57), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n658), .A2(KEYINPUT57), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n853), .B1(new_n852), .B2(new_n864), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n952), .B(new_n953), .C1(new_n875), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n656), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n771), .B(KEYINPUT122), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n939), .B1(new_n956), .B2(new_n958), .ZN(G54));
  INV_X1    g773(.A(KEYINPUT58), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n960), .A2(new_n348), .A3(KEYINPUT123), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n188), .B(new_n961), .C1(new_n852), .C2(new_n864), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT123), .B1(new_n960), .B2(new_n348), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n401), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n401), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n939), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(G60));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT59), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n617), .B1(new_n877), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n617), .B(new_n971), .C1(new_n875), .C2(new_n954), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n940), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n973), .B2(new_n940), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n852), .B2(new_n864), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n939), .B1(new_n980), .B2(new_n637), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n233), .B2(new_n980), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G66));
  NAND4_X1  g798(.A1(new_n830), .A2(new_n602), .A3(new_n642), .A4(new_n837), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n222), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n541), .B2(new_n570), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n946), .B1(G898), .B2(new_n222), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  OAI21_X1  g806(.A(G953), .B1(new_n516), .B2(new_n650), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n741), .A2(new_n812), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n779), .B1(new_n767), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n790), .A2(new_n854), .A3(new_n866), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n995), .A2(new_n996), .A3(new_n222), .A4(new_n751), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n317), .A2(new_n319), .ZN(new_n998));
  INV_X1    g812(.A(new_n390), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n203), .A2(KEYINPUT88), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT19), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n998), .B(new_n1003), .Z(new_n1004));
  NAND2_X1  g818(.A1(G900), .A2(G953), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n997), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n805), .A2(new_n672), .ZN(new_n1009));
  OR3_X1    g823(.A1(new_n696), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n696), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n676), .A2(new_n347), .A3(new_n763), .A4(new_n836), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n780), .A3(new_n790), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1004), .B1(new_n1014), .B2(new_n222), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n992), .B(new_n993), .C1(new_n1007), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1015), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n993), .A2(new_n992), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n993), .A2(new_n992), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1006), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1016), .A2(new_n1020), .ZN(G72));
  INV_X1    g835(.A(new_n343), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1014), .B2(new_n986), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n341), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n995), .A2(new_n996), .A3(new_n751), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1024), .B1(new_n1027), .B2(new_n986), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n342), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1022), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n343), .A2(new_n325), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n873), .A2(new_n1024), .A3(new_n1031), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n1030), .A2(new_n939), .A3(new_n1032), .ZN(G57));
endmodule


