//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT65), .ZN(new_n468));
  AND4_X1   g043(.A1(G137), .A2(new_n461), .A3(new_n463), .A4(new_n459), .ZN(new_n469));
  NOR3_X1   g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(G160));
  NAND3_X1  g045(.A1(new_n461), .A2(new_n463), .A3(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n461), .A2(new_n463), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n473), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n485), .A2(new_n461), .A3(new_n463), .A4(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n459), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n459), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G50), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT68), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n496), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(new_n497), .B2(new_n498), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G88), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n508), .B1(new_n503), .B2(new_n505), .ZN(new_n509));
  AND2_X1   g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n513), .B(G651), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n501), .B(new_n507), .C1(new_n512), .C2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND2_X1  g092(.A1(new_n506), .A2(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n499), .A2(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n503), .A2(new_n505), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n518), .A2(new_n520), .A3(new_n521), .A4(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  XOR2_X1   g100(.A(KEYINPUT71), .B(G90), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n506), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  INV_X1    g103(.A(new_n499), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n499), .A2(G43), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n497), .A2(new_n498), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n522), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n503), .B2(new_n505), .ZN(new_n550));
  AND2_X1   g125(.A1(G78), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g129(.A1(KEYINPUT6), .A2(G651), .ZN(new_n555));
  NOR2_X1   g130(.A1(KEYINPUT6), .A2(G651), .ZN(new_n556));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n558), .A2(new_n561), .B1(new_n506), .B2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  INV_X1    g138(.A(new_n561), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n557), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT73), .B(G651), .C1(new_n550), .C2(new_n551), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n554), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(G299));
  OAI221_X1 g142(.A(new_n527), .B1(new_n529), .B2(new_n528), .C1(new_n531), .C2(new_n532), .ZN(G301));
  AND3_X1   g143(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(G543), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n532), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT74), .B1(new_n539), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n506), .A2(new_n576), .A3(G87), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n499), .A2(G49), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G288));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n555), .C2(new_n556), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT77), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n538), .A2(new_n585), .A3(G48), .A4(G543), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n584), .B(new_n586), .C1(new_n539), .C2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n503), .B2(new_n505), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT76), .B(G651), .C1(new_n590), .C2(new_n592), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n588), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n532), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n499), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n539), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT10), .B1(new_n539), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n499), .A2(G54), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n503), .B2(new_n505), .ZN(new_n611));
  AND2_X1   g186(.A1(G79), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n506), .A2(new_n614), .A3(G92), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n608), .A2(new_n609), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G299), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  INV_X1    g200(.A(new_n542), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n620), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n475), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n472), .A2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n462), .A2(new_n460), .A3(G2105), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT13), .B(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n636), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(G14), .ZN(G401));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT81), .Z(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT17), .Z(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT80), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT82), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n657), .A3(new_n659), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  INV_X1    g241(.A(new_n659), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n658), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n662), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n668), .B(new_n669), .C1(new_n658), .C2(new_n660), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2100), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n676), .A2(new_n679), .A3(new_n681), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(new_n683), .C2(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT22), .B(G1981), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n688), .A2(new_n690), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n701));
  INV_X1    g276(.A(G26), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G29), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n475), .A2(G140), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  INV_X1    g281(.A(G128), .ZN(new_n707));
  NOR2_X1   g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n471), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n704), .B1(new_n711), .B2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n703), .B1(new_n712), .B2(new_n701), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(G2067), .ZN(new_n714));
  INV_X1    g289(.A(G11), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(G2067), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n714), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G168), .A2(G16), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n720), .B1(new_n721), .B2(G1966), .C1(G16), .C2(G21), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(G1966), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G171), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G5), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n475), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n472), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  NAND4_X1  g307(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G29), .B2(G32), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n726), .A2(new_n727), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G34), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(G34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n742), .A2(new_n743), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G160), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n738), .B1(new_n727), .B2(new_n726), .C1(new_n739), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(G299), .A2(G16), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n752), .A2(KEYINPUT23), .A3(G20), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n754));
  INV_X1    g329(.A(G20), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G16), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n635), .A2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT95), .B(G28), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT30), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n761), .B1(new_n740), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n749), .A2(new_n739), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n759), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n719), .A2(new_n724), .A3(new_n750), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n752), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n617), .B2(new_n752), .ZN(new_n769));
  INV_X1    g344(.A(G1348), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G164), .A2(new_n740), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G27), .B2(new_n740), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(new_n736), .B2(new_n737), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n767), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G29), .B2(G33), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n778), .A2(G29), .A3(G33), .ZN(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G127), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n474), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2105), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT25), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n475), .A2(G139), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n779), .B(new_n780), .C1(new_n788), .C2(new_n740), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2072), .Z(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n740), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n740), .ZN(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n752), .A2(G19), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n542), .B2(new_n752), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1341), .Z(new_n800));
  NAND4_X1  g375(.A1(new_n777), .A2(new_n791), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n802));
  NAND2_X1  g377(.A1(G288), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT87), .A3(new_n581), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n752), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT33), .B(G1976), .Z(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G23), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n752), .A2(G22), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G303), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1971), .ZN(new_n814));
  INV_X1    g389(.A(new_n807), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n805), .B2(new_n808), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n752), .A2(G6), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n597), .B2(new_n752), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT32), .B(G1981), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n810), .A2(new_n814), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n475), .A2(G131), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n826));
  INV_X1    g401(.A(G95), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n459), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT84), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n459), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(KEYINPUT84), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n825), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G119), .ZN(new_n835));
  OR3_X1    g410(.A1(new_n471), .A2(KEYINPUT83), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT83), .B1(new_n471), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT85), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n828), .A2(new_n829), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n832), .A2(KEYINPUT84), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n840), .A2(new_n841), .B1(G131), .B2(new_n475), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT85), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n837), .A4(new_n836), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT86), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT86), .B1(new_n839), .B2(new_n844), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n847), .A2(new_n740), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(G25), .A2(G29), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n824), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n824), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n845), .B(new_n846), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n740), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n752), .A2(G24), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n604), .B2(new_n752), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(G1986), .Z(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n859), .C1(new_n821), .C2(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT88), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n810), .A2(new_n816), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT34), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n814), .A4(new_n820), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT88), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n859), .A4(new_n856), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n823), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT89), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(KEYINPUT36), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(KEYINPUT36), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n801), .B1(new_n871), .B2(new_n872), .ZN(G311));
  NOR2_X1   g448(.A1(new_n867), .A2(new_n870), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n869), .B(new_n823), .C1(new_n861), .C2(new_n866), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n777), .A2(new_n800), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n876), .A2(new_n791), .A3(new_n797), .A4(new_n877), .ZN(G150));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n522), .A2(G67), .ZN(new_n880));
  AND2_X1   g455(.A1(G80), .A2(G543), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n879), .B(G651), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n522), .B2(G67), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT97), .B1(new_n883), .B2(new_n532), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT98), .B(G55), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n499), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G93), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n539), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(KEYINPUT99), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(KEYINPUT99), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT100), .B(G860), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT37), .Z(new_n895));
  NOR2_X1   g470(.A1(new_n892), .A2(new_n542), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n889), .B(KEYINPUT99), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n626), .B1(new_n897), .B2(new_n885), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n616), .A2(new_n624), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n895), .B1(new_n903), .B2(new_n893), .ZN(G145));
  INV_X1    g479(.A(new_n635), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n480), .A2(new_n748), .A3(new_n481), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n748), .B1(new_n480), .B2(new_n481), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n635), .A3(new_n906), .ZN(new_n911));
  INV_X1    g486(.A(new_n639), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n909), .B2(new_n911), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n845), .A2(new_n734), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n839), .A2(new_n844), .A3(new_n733), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n484), .A2(KEYINPUT4), .A3(G138), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n487), .B1(new_n474), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n459), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n492), .A2(new_n493), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G2105), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n489), .A2(new_n490), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n919), .A2(new_n926), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n459), .A2(G118), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT102), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n475), .A2(G142), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n472), .A2(G130), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n928), .A2(new_n929), .A3(new_n936), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G164), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n939), .B2(new_n927), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n918), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n936), .B1(new_n928), .B2(new_n929), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n927), .A3(new_n935), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n917), .A3(new_n916), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n944), .A3(new_n711), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n711), .B1(new_n941), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n915), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n944), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n706), .A2(new_n710), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n951), .B(new_n945), .C1(new_n914), .C2(new_n913), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g530(.A(new_n899), .B(new_n628), .ZN(new_n956));
  NAND2_X1  g531(.A1(G299), .A2(KEYINPUT103), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n558), .A2(new_n561), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n506), .A2(G91), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n958), .A2(new_n565), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n554), .A4(new_n566), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n962), .A3(new_n616), .ZN(new_n963));
  OR3_X1    g538(.A1(G299), .A2(KEYINPUT103), .A3(new_n616), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n956), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(KEYINPUT41), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n964), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n956), .A2(new_n967), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(new_n973), .B2(KEYINPUT104), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n966), .A2(KEYINPUT104), .ZN(new_n975));
  AOI21_X1  g550(.A(G290), .B1(new_n803), .B2(new_n804), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n803), .A2(G290), .A3(new_n804), .ZN(new_n978));
  AOI21_X1  g553(.A(G305), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n978), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n980), .A2(new_n976), .A3(new_n597), .ZN(new_n981));
  OAI21_X1  g556(.A(G303), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n597), .B1(new_n980), .B2(new_n976), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(G305), .A3(new_n978), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(G166), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n988));
  AND4_X1   g563(.A1(new_n974), .A2(new_n975), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n975), .A2(new_n974), .B1(new_n987), .B2(new_n988), .ZN(new_n990));
  OAI21_X1  g565(.A(G868), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n892), .A2(new_n620), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(G295));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n992), .ZN(G331));
  XOR2_X1   g569(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n995));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n996));
  NAND2_X1  g571(.A1(G171), .A2(G286), .ZN(new_n997));
  NAND2_X1  g572(.A1(G168), .A2(G301), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n896), .A2(new_n898), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n892), .A2(new_n542), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n897), .A2(new_n626), .A3(new_n885), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n1001), .A2(new_n1002), .B1(new_n998), .B2(new_n997), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n996), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n999), .B1(new_n896), .B2(new_n898), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT107), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1004), .A2(new_n964), .A3(new_n963), .A4(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1001), .A2(new_n1002), .A3(new_n998), .A4(new_n997), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n972), .A2(new_n967), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n982), .A3(new_n1010), .A4(new_n985), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n953), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1010), .A2(new_n1007), .B1(new_n982), .B2(new_n985), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n995), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1004), .A2(new_n1006), .B1(new_n968), .B2(new_n971), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1009), .A2(new_n965), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n986), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n995), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1011), .A3(new_n953), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(KEYINPUT44), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1012), .A2(new_n1013), .A3(new_n995), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1011), .A3(new_n953), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(KEYINPUT44), .B2(new_n1025), .ZN(G397));
  NOR2_X1   g601(.A1(new_n845), .A2(new_n853), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT108), .B(G1384), .Z(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n926), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G40), .ZN(new_n1030));
  NOR4_X1   g605(.A1(new_n466), .A2(new_n468), .A3(new_n1030), .A4(new_n469), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n824), .B1(new_n839), .B2(new_n844), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1027), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1996), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n734), .ZN(new_n1039));
  INV_X1    g614(.A(G2067), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n950), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(G1996), .B2(new_n733), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n711), .A2(G2067), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1039), .B1(new_n1033), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n604), .B(G1986), .Z(new_n1047));
  AOI211_X1 g622(.A(new_n1035), .B(new_n1046), .C1(new_n1032), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1384), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n926), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G160), .A2(G40), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT113), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1031), .A2(new_n1049), .A3(new_n926), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT118), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n506), .A2(G86), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1060), .A2(new_n584), .A3(new_n586), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1061), .B2(new_n593), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT115), .B(G1981), .Z(new_n1064));
  OAI21_X1  g639(.A(G61), .B1(new_n569), .B2(new_n570), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n591), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT76), .B1(new_n1066), .B2(G651), .ZN(new_n1067));
  INV_X1    g642(.A(new_n596), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1061), .B(new_n1064), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n597), .B2(new_n1064), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1063), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n597), .A2(KEYINPUT116), .A3(new_n1064), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1063), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(new_n1057), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G288), .A2(G1976), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1081), .B(KEYINPUT119), .Z(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1058), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n803), .A2(new_n804), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1057), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT49), .B1(new_n1078), .B2(new_n1063), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1074), .B(new_n1062), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1091), .B2(new_n1057), .ZN(new_n1092));
  INV_X1    g667(.A(G1971), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n926), .A2(KEYINPUT45), .A3(new_n1028), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1031), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT45), .B1(new_n926), .B2(new_n1049), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT110), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1050), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n926), .A2(KEYINPUT50), .A3(new_n1049), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1051), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n794), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n926), .A2(KEYINPUT50), .A3(new_n1049), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT50), .B1(new_n926), .B2(new_n1049), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n794), .B(new_n1031), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT111), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(new_n1093), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1098), .A2(new_n1104), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT55), .ZN(new_n1115));
  INV_X1    g690(.A(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(G166), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1111), .A2(G8), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1097), .B2(new_n1107), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT114), .B(G1976), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT52), .B1(G288), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1057), .A2(new_n1087), .A3(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1092), .A2(new_n1120), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(G299), .B(KEYINPUT57), .Z(new_n1127));
  OAI21_X1  g702(.A(new_n1031), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n758), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT45), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(G164), .B2(G1384), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT56), .B(G2072), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1031), .A3(new_n1094), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT123), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1127), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1050), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1040), .A4(new_n1031), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1031), .A2(new_n1049), .A3(new_n1040), .A4(new_n926), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(new_n770), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1129), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1148), .A2(new_n617), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1139), .A2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n616), .B(KEYINPUT124), .Z(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1147), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1102), .A2(G1348), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1145), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1155), .A2(new_n1145), .A3(new_n1154), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n616), .A2(KEYINPUT124), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1153), .B(new_n1156), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1131), .A2(new_n1036), .A3(new_n1031), .A4(new_n1094), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1054), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT58), .B(G1341), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n542), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(new_n1166), .A3(new_n542), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1127), .B1(new_n1133), .B2(new_n1129), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1149), .B1(new_n1169), .B2(KEYINPUT61), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1135), .A2(new_n1171), .A3(new_n1127), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1159), .A2(new_n1168), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1126), .B1(new_n1151), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT51), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(KEYINPUT125), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G286), .A2(G8), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT120), .B(G2084), .Z(new_n1179));
  NAND3_X1  g754(.A1(new_n926), .A2(KEYINPUT45), .A3(new_n1049), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1131), .A2(new_n1031), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(G1966), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1102), .A2(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1177), .B(new_n1178), .C1(new_n1183), .C2(new_n1116), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1031), .B(new_n1179), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n926), .A2(KEYINPUT45), .A3(new_n1049), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1186), .A2(new_n1096), .A3(new_n1051), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1185), .B1(new_n1187), .B2(G1966), .ZN(new_n1188));
  OAI211_X1 g763(.A(G8), .B(new_n1176), .C1(new_n1188), .C2(G286), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1175), .A2(KEYINPUT125), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1184), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1183), .A2(new_n1116), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(G286), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1187), .A2(KEYINPUT53), .A3(new_n774), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT53), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1131), .A2(new_n1031), .A3(new_n1094), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(G2078), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1128), .A2(new_n727), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(G301), .B(KEYINPUT54), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OR4_X1    g777(.A1(new_n1196), .A2(new_n1095), .A3(G2078), .A4(new_n1029), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1201), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1203), .A2(new_n1198), .A3(new_n1199), .A4(new_n1204), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1194), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1084), .B1(new_n1174), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1194), .A2(KEYINPUT62), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(KEYINPUT126), .ZN(new_n1209));
  OR2_X1    g784(.A1(new_n1194), .A2(KEYINPUT62), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1194), .A2(new_n1211), .A3(KEYINPUT62), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1200), .A2(G171), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1126), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1057), .A2(new_n1087), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(KEYINPUT52), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1080), .A2(new_n1217), .A3(new_n1125), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(KEYINPUT117), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT117), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1080), .A2(new_n1217), .A3(new_n1220), .A4(new_n1125), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  OR2_X1    g797(.A1(new_n1222), .A2(new_n1120), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1207), .A2(new_n1215), .A3(new_n1223), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1080), .A2(new_n1217), .A3(new_n1125), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1192), .A2(G168), .ZN(new_n1226));
  INV_X1    g801(.A(new_n1226), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1225), .A2(new_n1120), .A3(new_n1122), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT121), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT63), .ZN(new_n1230));
  AND3_X1   g805(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1111), .A2(G8), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1119), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1234), .A2(KEYINPUT63), .A3(new_n1120), .ZN(new_n1235));
  NOR3_X1   g810(.A1(new_n1222), .A2(new_n1235), .A3(new_n1226), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1229), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1237));
  NOR3_X1   g812(.A1(new_n1231), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1048), .B1(new_n1224), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g814(.A(KEYINPUT46), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n1038), .B(new_n1240), .ZN(new_n1241));
  AND3_X1   g816(.A1(new_n1044), .A2(new_n734), .A3(new_n1041), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1241), .B1(new_n1033), .B2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT47), .ZN(new_n1244));
  NOR3_X1   g819(.A1(new_n1046), .A2(new_n854), .A3(new_n824), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1032), .B1(new_n1245), .B2(new_n1042), .ZN(new_n1246));
  NOR3_X1   g821(.A1(new_n1033), .A2(G1986), .A3(G290), .ZN(new_n1247));
  XNOR2_X1  g822(.A(new_n1247), .B(KEYINPUT48), .ZN(new_n1248));
  OR3_X1    g823(.A1(new_n1046), .A2(new_n1035), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g824(.A1(new_n1244), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g825(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1239), .A2(new_n1251), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g827(.A1(new_n954), .A2(new_n699), .A3(new_n673), .ZN(new_n1254));
  INV_X1    g828(.A(G319), .ZN(new_n1255));
  AOI21_X1  g829(.A(new_n1255), .B1(new_n655), .B2(G14), .ZN(new_n1256));
  NAND3_X1  g830(.A1(new_n1020), .A2(new_n1254), .A3(new_n1256), .ZN(G225));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1258));
  NAND2_X1  g832(.A1(G225), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g833(.A1(new_n1020), .A2(new_n1254), .A3(KEYINPUT127), .A4(new_n1256), .ZN(new_n1260));
  NAND2_X1  g834(.A1(new_n1259), .A2(new_n1260), .ZN(G308));
endmodule


