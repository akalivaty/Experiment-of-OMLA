//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G101), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G137), .A3(new_n461), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n461), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n475), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n480), .B2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n480), .A2(new_n461), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n465), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n487), .A2(G124), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n473), .A2(new_n475), .A3(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n466), .A2(G102), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT68), .A2(G138), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n473), .A2(new_n475), .A3(new_n499), .A4(new_n461), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n470), .A2(KEYINPUT4), .A3(new_n461), .A4(new_n499), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(new_n498), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT69), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n511), .A2(G50), .A3(G543), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n508), .A2(new_n510), .B1(KEYINPUT6), .B2(new_n507), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .A3(G50), .A4(G543), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n515), .A2(new_n517), .B1(new_n524), .B2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(KEYINPUT71), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND3_X1  g110(.A1(new_n516), .A2(G89), .A3(new_n523), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n511), .A2(G543), .A3(new_n512), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G51), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n538), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n538), .A2(new_n543), .A3(new_n546), .A4(new_n540), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n524), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n542), .A2(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n522), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(new_n524), .A2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n542), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n522), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT73), .ZN(G188));
  NAND4_X1  g146(.A1(new_n511), .A2(G53), .A3(G543), .A4(new_n512), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n524), .A2(G91), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n522), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(G299));
  AND2_X1   g156(.A1(new_n545), .A2(new_n547), .ZN(G286));
  NAND3_X1  g157(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n516), .A2(G87), .A3(new_n523), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT74), .Z(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n522), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n516), .A2(G86), .A3(new_n523), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n522), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT75), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n524), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n542), .A2(G47), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n516), .A2(new_n523), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n522), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n605), .A2(new_n609), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n542), .A2(G54), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G284));
  XNOR2_X1  g191(.A(G284), .B(KEYINPUT76), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g202(.A1(new_n480), .A2(new_n462), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  NAND2_X1  g206(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n636), .B(new_n637), .C1(G111), .C2(new_n461), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n487), .A2(G123), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n482), .A2(new_n484), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  OAI211_X1 g219(.A(new_n633), .B(new_n644), .C1(KEYINPUT78), .C2(G2100), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2443), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT17), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n669), .C2(new_n665), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n682), .B1(KEYINPUT20), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(KEYINPUT20), .C2(new_n684), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT83), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(G229));
  AND3_X1   g269(.A1(G168), .A2(KEYINPUT91), .A3(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT91), .B1(G168), .B2(G16), .ZN(new_n696));
  OAI22_X1  g271(.A1(new_n695), .A2(new_n696), .B1(G16), .B2(G21), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1966), .ZN(new_n698));
  AND2_X1   g273(.A1(KEYINPUT84), .A2(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(KEYINPUT84), .A2(G29), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G299), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT23), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G20), .ZN(new_n711));
  MUX2_X1   g286(.A(KEYINPUT23), .B(new_n710), .S(new_n711), .Z(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(G1956), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n705), .A2(new_n706), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n707), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(G29), .A2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n487), .A2(G129), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n485), .A2(G141), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n466), .A2(G105), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n719), .A2(new_n720), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n716), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT27), .B(G1996), .ZN(new_n727));
  NOR2_X1   g302(.A1(G5), .A2(G16), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G171), .B2(G16), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n726), .A2(new_n727), .B1(G1961), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n701), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n701), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G34), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n701), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G160), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n725), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(G28), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT30), .B2(new_n744), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n643), .B2(new_n701), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n730), .A2(new_n734), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n709), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n615), .B2(new_n709), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1348), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n749), .B(new_n752), .C1(G1956), .C2(new_n712), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n729), .A2(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n701), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n485), .A2(G140), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  INV_X1    g334(.A(G116), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n465), .B1(new_n760), .B2(G2105), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n487), .A2(G128), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(new_n725), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g342(.A(G2067), .B(new_n757), .C1(new_n764), .C2(new_n725), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n754), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n725), .A2(G33), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n482), .A2(G139), .A3(new_n484), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n466), .A2(G103), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT89), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n771), .A2(new_n776), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  INV_X1    g353(.A(G127), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n480), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n775), .A2(new_n777), .B1(G2105), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n770), .B1(new_n781), .B2(new_n725), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G2072), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n769), .B(new_n783), .C1(new_n726), .C2(new_n727), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n709), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n564), .B2(new_n709), .ZN(new_n786));
  MUX2_X1   g361(.A(new_n785), .B(new_n786), .S(KEYINPUT87), .Z(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G1341), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(G1341), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n782), .B2(G2072), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n784), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AND4_X1   g367(.A1(new_n698), .A2(new_n715), .A3(new_n753), .A4(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT31), .B(G11), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n709), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(new_n586), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n709), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(KEYINPUT33), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(KEYINPUT33), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n801), .A2(G1976), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(G1976), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n709), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n709), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G1971), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(G1971), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n709), .A2(G6), .ZN(new_n810));
  INV_X1    g385(.A(G305), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n709), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT86), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n808), .A2(new_n809), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n796), .B1(new_n805), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n808), .A2(new_n809), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n803), .A2(new_n804), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT34), .A4(new_n815), .ZN(new_n820));
  AND2_X1   g395(.A1(G290), .A2(KEYINPUT85), .ZN(new_n821));
  NOR2_X1   g396(.A1(G290), .A2(KEYINPUT85), .ZN(new_n822));
  OAI21_X1  g397(.A(G16), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G16), .B2(G24), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(G1986), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(G1986), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n817), .A2(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  OR2_X1    g403(.A1(G95), .A2(G2105), .ZN(new_n829));
  INV_X1    g404(.A(G107), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n465), .B1(new_n830), .B2(G2105), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n487), .A2(G119), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G131), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n642), .B2(new_n833), .ZN(new_n834));
  MUX2_X1   g409(.A(new_n834), .B(G25), .S(new_n701), .Z(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT35), .B(G1991), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n827), .A2(new_n828), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n828), .B1(new_n827), .B2(new_n838), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n793), .B(new_n795), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT93), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n827), .A2(new_n838), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n827), .A2(new_n828), .A3(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n847), .A2(new_n848), .A3(new_n795), .A4(new_n793), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n843), .A2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n522), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G651), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI221_X1 g431(.A(new_n854), .B1(new_n855), .B2(new_n541), .C1(new_n856), .C2(new_n607), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n613), .A2(new_n614), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n622), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(KEYINPUT94), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n542), .A2(G55), .B1(G651), .B2(new_n853), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n865), .B(new_n866), .C1(new_n856), .C2(new_n607), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n867), .A3(new_n564), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n564), .B1(new_n864), .B2(new_n867), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n863), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n859), .B1(new_n872), .B2(G860), .ZN(G145));
  OR2_X1    g448(.A1(new_n461), .A2(G118), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n465), .B1(new_n874), .B2(KEYINPUT97), .ZN(new_n875));
  OAI221_X1 g450(.A(new_n875), .B1(KEYINPUT97), .B2(new_n874), .C1(G106), .C2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(G130), .ZN(new_n877));
  INV_X1    g452(.A(new_n487), .ZN(new_n878));
  INV_X1    g453(.A(G142), .ZN(new_n879));
  OAI221_X1 g454(.A(new_n876), .B1(new_n877), .B2(new_n878), .C1(new_n642), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n834), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(new_n630), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n630), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(KEYINPUT98), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n881), .A2(new_n630), .ZN(new_n886));
  INV_X1    g461(.A(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n834), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n880), .B(new_n832), .C1(new_n833), .C2(new_n642), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(new_n630), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n885), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n775), .A2(new_n777), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n780), .A2(G2105), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(KEYINPUT96), .A3(new_n763), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n764), .B1(new_n781), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n898), .A3(new_n724), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n724), .B1(new_n896), .B2(new_n898), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n504), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n898), .ZN(new_n903));
  INV_X1    g478(.A(new_n724), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G164), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n892), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n504), .B1(new_n900), .B2(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n884), .A2(new_n891), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(G164), .A3(new_n899), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(KEYINPUT99), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n492), .B(KEYINPUT95), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n915), .A2(G160), .ZN(new_n916));
  INV_X1    g491(.A(new_n643), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(G160), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n908), .A2(new_n910), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n892), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n908), .A2(new_n910), .A3(new_n883), .A4(new_n882), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g503(.A1(new_n857), .A2(new_n618), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n624), .B(KEYINPUT100), .Z(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n871), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n624), .B(KEYINPUT100), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n869), .B2(new_n870), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n615), .A2(new_n708), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n860), .A2(G299), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n932), .B(new_n871), .ZN(new_n938));
  INV_X1    g513(.A(new_n935), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n860), .A2(G299), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT41), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n937), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G290), .A2(new_n798), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(G290), .A2(new_n798), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(G166), .ZN(new_n949));
  OR2_X1    g524(.A1(G290), .A2(new_n798), .ZN(new_n950));
  AOI21_X1  g525(.A(G303), .B1(new_n950), .B2(new_n946), .ZN(new_n951));
  OAI21_X1  g526(.A(G305), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(G166), .B1(new_n947), .B2(new_n948), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n946), .A3(G303), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n811), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(KEYINPUT101), .A3(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n957), .A2(KEYINPUT101), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(KEYINPUT101), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n952), .A2(new_n955), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n945), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n929), .B1(new_n963), .B2(new_n618), .ZN(G295));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(new_n929), .C1(new_n963), .C2(new_n618), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n945), .A2(new_n961), .A3(new_n958), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n931), .A2(new_n933), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n943), .A3(new_n941), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n969), .A3(new_n937), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n618), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n929), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT102), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(G331));
  INV_X1    g549(.A(new_n936), .ZN(new_n975));
  OAI21_X1  g550(.A(G286), .B1(new_n869), .B2(new_n870), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n864), .A2(new_n867), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n563), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(G168), .A3(new_n868), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n976), .A2(new_n979), .A3(G171), .ZN(new_n980));
  AOI21_X1  g555(.A(G171), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n869), .A2(G286), .A3(new_n870), .ZN(new_n983));
  AOI21_X1  g558(.A(G168), .B1(new_n978), .B2(new_n868), .ZN(new_n984));
  OAI21_X1  g559(.A(G301), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n976), .A2(new_n979), .A3(G171), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n944), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n987), .A3(new_n956), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n982), .A2(new_n987), .A3(new_n956), .A4(KEYINPUT105), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G37), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n982), .A2(new_n987), .ZN(new_n995));
  INV_X1    g570(.A(new_n956), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n941), .A2(KEYINPUT106), .A3(new_n943), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n936), .A2(new_n1000), .A3(KEYINPUT41), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n985), .A2(new_n999), .A3(new_n986), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n982), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n996), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n990), .A2(new_n1004), .A3(new_n993), .A4(new_n991), .ZN(new_n1005));
  INV_X1    g580(.A(new_n994), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n998), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n990), .A2(new_n997), .A3(new_n993), .A4(new_n991), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1010), .B(KEYINPUT44), .C1(new_n994), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(G397));
  NAND4_X1  g588(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(G1976), .ZN(new_n1014));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  INV_X1    g590(.A(new_n495), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n470), .B2(G126), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n498), .B1(new_n1017), .B2(new_n461), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n502), .A2(new_n503), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n478), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT107), .B(G40), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1021), .A2(new_n471), .A3(new_n469), .A4(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1014), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT112), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n472), .A2(new_n478), .A3(new_n1022), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1015), .A3(new_n504), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(G8), .A4(new_n1014), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1030), .A3(KEYINPUT52), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n592), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1034), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1028), .A2(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1037), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1025), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1045), .B(new_n1046), .C1(new_n587), .C2(G1976), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1026), .A2(new_n1030), .A3(KEYINPUT113), .A4(KEYINPUT52), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1033), .A2(new_n1044), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1043), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(KEYINPUT115), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n1015), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n504), .B2(new_n1015), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(KEYINPUT110), .A3(new_n706), .A4(new_n1027), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1020), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1027), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1971), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(new_n706), .A3(new_n1027), .A4(new_n1055), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1059), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1071), .B(new_n1072), .C1(G166), .C2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n525), .B2(new_n533), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT55), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT111), .B1(new_n1075), .B2(KEYINPUT55), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1070), .A2(new_n1078), .A3(G8), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1051), .A2(new_n1053), .A3(new_n1079), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1043), .A2(G1976), .A3(G288), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G305), .A2(G1981), .ZN(new_n1082));
  OAI211_X1 g657(.A(G8), .B(new_n1028), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1073), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1079), .A2(new_n1049), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  INV_X1    g663(.A(G1966), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1063), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1066), .A2(new_n741), .A3(new_n1027), .A4(new_n1055), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1092), .B2(G286), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(G168), .A3(new_n1091), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1088), .B1(new_n1094), .B2(G8), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT62), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1061), .A2(new_n733), .A3(new_n1027), .A4(new_n1062), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1066), .A2(new_n1027), .A3(new_n1055), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1100), .A2(G2078), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1061), .A2(new_n1027), .A3(new_n1062), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1095), .A2(KEYINPUT51), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1109), .B(new_n1110), .C1(new_n1095), .C2(new_n1093), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1087), .A2(new_n1098), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT124), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1108), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1092), .A2(G286), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1094), .A2(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1097), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1114), .B1(new_n1118), .B2(new_n1110), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1087), .A4(new_n1098), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1084), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1117), .A2(G168), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1117), .B2(G168), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G299), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n575), .A2(KEYINPUT57), .A3(new_n576), .A4(new_n580), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT120), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1102), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1061), .A2(new_n1027), .A3(new_n1062), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1027), .A2(KEYINPUT118), .A3(new_n1015), .A4(new_n504), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n766), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1348), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1102), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT119), .A4(new_n766), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n615), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(KEYINPUT121), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1138), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1153), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .A4(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(G1996), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1160), .A2(new_n1061), .A3(new_n1027), .A4(new_n1062), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT58), .B(G1341), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n564), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT59), .B(new_n564), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1151), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1170), .A2(new_n860), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1149), .B(new_n615), .C1(new_n1150), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n860), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1139), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n1177));
  INV_X1    g752(.A(G40), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n476), .A2(new_n477), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT122), .Z(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1180), .B2(G2105), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n472), .A2(new_n1100), .A3(G2078), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1061), .A3(new_n1062), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1101), .A2(new_n1104), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1184), .A2(G171), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1177), .B1(new_n1108), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1109), .B1(new_n1095), .B2(new_n1093), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1184), .A2(G171), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1101), .A2(new_n1104), .A3(G301), .A4(new_n1107), .ZN(new_n1190));
  AND4_X1   g765(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT54), .A4(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1177), .B1(new_n1184), .B2(G171), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1188), .B1(new_n1192), .B2(new_n1190), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1186), .B(new_n1187), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1128), .B1(new_n1176), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1087), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1070), .A2(G8), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1078), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1051), .A2(new_n1053), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT117), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1124), .B(KEYINPUT116), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1051), .A2(new_n1053), .A3(KEYINPUT117), .A4(new_n1199), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1079), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(KEYINPUT63), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1122), .A2(new_n1196), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n724), .B(new_n1160), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n763), .B(new_n766), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n834), .B(new_n837), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1061), .A2(new_n1024), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(G290), .A2(G1986), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT108), .Z(new_n1217));
  AOI21_X1  g792(.A(new_n1217), .B1(G1986), .B2(G290), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1214), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1215), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT109), .Z(new_n1221));
  NAND2_X1  g796(.A1(new_n1208), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1214), .A2(new_n1160), .ZN(new_n1223));
  XOR2_X1   g798(.A(new_n1223), .B(KEYINPUT46), .Z(new_n1224));
  AOI21_X1  g799(.A(new_n1219), .B1(new_n1210), .B2(new_n904), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1226), .B(new_n1227), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n834), .A2(new_n836), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1211), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n764), .A2(new_n766), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1219), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n1233));
  XNOR2_X1  g808(.A(new_n1232), .B(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1217), .A2(new_n1214), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n1235), .B(KEYINPUT48), .ZN(new_n1236));
  AOI211_X1 g811(.A(new_n1228), .B(new_n1234), .C1(new_n1215), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1222), .A2(new_n1237), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g813(.A(G319), .ZN(new_n1240));
  OR3_X1    g814(.A1(G229), .A2(new_n1240), .A3(G227), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1241), .B1(new_n922), .B2(new_n926), .ZN(new_n1242));
  AND4_X1   g816(.A1(new_n660), .A2(new_n1242), .A3(new_n998), .A4(new_n1007), .ZN(G308));
  NAND4_X1  g817(.A1(new_n1242), .A2(new_n998), .A3(new_n660), .A4(new_n1007), .ZN(G225));
endmodule


