

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582;

  INV_X1 U319 ( .A(KEYINPUT108), .ZN(n399) );
  XNOR2_X1 U320 ( .A(n305), .B(n304), .ZN(n332) );
  XNOR2_X1 U321 ( .A(n459), .B(n458), .ZN(n513) );
  XNOR2_X1 U322 ( .A(n457), .B(KEYINPUT93), .ZN(n458) );
  XNOR2_X1 U323 ( .A(n437), .B(KEYINPUT109), .ZN(n529) );
  XOR2_X1 U324 ( .A(n550), .B(KEYINPUT28), .Z(n520) );
  XOR2_X1 U325 ( .A(n308), .B(n307), .Z(n287) );
  INV_X1 U326 ( .A(KEYINPUT106), .ZN(n355) );
  INV_X1 U327 ( .A(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U328 ( .A(n303), .B(n302), .ZN(n305) );
  INV_X1 U329 ( .A(KEYINPUT37), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n405), .B(n404), .ZN(n411) );
  XNOR2_X1 U331 ( .A(n411), .B(n410), .ZN(n415) );
  XNOR2_X1 U332 ( .A(n317), .B(KEYINPUT36), .ZN(n318) );
  XNOR2_X1 U333 ( .A(n309), .B(n287), .ZN(n310) );
  XNOR2_X1 U334 ( .A(n567), .B(n318), .ZN(n578) );
  XNOR2_X1 U335 ( .A(n311), .B(n310), .ZN(n316) );
  INV_X1 U336 ( .A(G127GAT), .ZN(n439) );
  XOR2_X1 U337 ( .A(n434), .B(n433), .Z(n554) );
  XNOR2_X1 U338 ( .A(n439), .B(KEYINPUT50), .ZN(n440) );
  XNOR2_X1 U339 ( .A(n463), .B(G43GAT), .ZN(n464) );
  XNOR2_X1 U340 ( .A(n441), .B(n440), .ZN(G1342GAT) );
  XNOR2_X1 U341 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT74), .B(G64GAT), .Z(n289) );
  XNOR2_X1 U343 ( .A(G127GAT), .B(G211GAT), .ZN(n288) );
  XNOR2_X1 U344 ( .A(n289), .B(n288), .ZN(n292) );
  XNOR2_X1 U345 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n290) );
  XNOR2_X1 U346 ( .A(n290), .B(KEYINPUT12), .ZN(n291) );
  XOR2_X1 U347 ( .A(n292), .B(n291), .Z(n294) );
  NAND2_X1 U348 ( .A1(G231GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n301) );
  XOR2_X1 U350 ( .A(G8GAT), .B(G183GAT), .Z(n366) );
  XOR2_X1 U351 ( .A(KEYINPUT13), .B(G57GAT), .Z(n296) );
  XNOR2_X1 U352 ( .A(G71GAT), .B(G78GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n340) );
  XOR2_X1 U354 ( .A(n366), .B(n340), .Z(n299) );
  XNOR2_X1 U355 ( .A(G15GAT), .B(G1GAT), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n297), .B(KEYINPUT66), .ZN(n328) );
  XOR2_X1 U357 ( .A(G22GAT), .B(G155GAT), .Z(n406) );
  XNOR2_X1 U358 ( .A(n328), .B(n406), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n479) );
  INV_X1 U361 ( .A(n479), .ZN(n575) );
  XOR2_X1 U362 ( .A(KEYINPUT104), .B(n575), .Z(n565) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(G29GAT), .ZN(n303) );
  XOR2_X1 U364 ( .A(KEYINPUT65), .B(KEYINPUT8), .Z(n304) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U366 ( .A(n332), .B(n404), .ZN(n311) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n306), .B(G218GAT), .ZN(n370) );
  XOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .Z(n341) );
  XOR2_X1 U370 ( .A(n370), .B(n341), .Z(n309) );
  XOR2_X1 U371 ( .A(G92GAT), .B(KEYINPUT9), .Z(n308) );
  NAND2_X1 U372 ( .A1(G232GAT), .A2(G233GAT), .ZN(n307) );
  XOR2_X1 U373 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n313) );
  XNOR2_X1 U374 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(n314), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n567) );
  INV_X1 U378 ( .A(KEYINPUT92), .ZN(n317) );
  OR2_X1 U379 ( .A1(n479), .A2(n578), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n319), .B(KEYINPUT45), .ZN(n354) );
  XOR2_X1 U381 ( .A(KEYINPUT64), .B(KEYINPUT68), .Z(n321) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n336) );
  XOR2_X1 U384 ( .A(G113GAT), .B(G50GAT), .Z(n323) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(G36GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U387 ( .A(KEYINPUT30), .B(G141GAT), .Z(n325) );
  XNOR2_X1 U388 ( .A(G22GAT), .B(G197GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U390 ( .A(n327), .B(n326), .Z(n334) );
  XOR2_X1 U391 ( .A(n328), .B(KEYINPUT67), .Z(n330) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n556) );
  INV_X1 U397 ( .A(n556), .ZN(n500) );
  XOR2_X1 U398 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n338) );
  XNOR2_X1 U399 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U401 ( .A(n340), .B(n339), .Z(n343) );
  XOR2_X1 U402 ( .A(G106GAT), .B(G148GAT), .Z(n407) );
  XNOR2_X1 U403 ( .A(n407), .B(n341), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U405 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n345) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(n347), .B(n346), .Z(n352) );
  XOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT71), .Z(n349) );
  XNOR2_X1 U410 ( .A(G176GAT), .B(G92GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U412 ( .A(G204GAT), .B(n350), .Z(n367) );
  XNOR2_X1 U413 ( .A(n367), .B(KEYINPUT32), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n572) );
  NAND2_X1 U415 ( .A1(n500), .A2(n572), .ZN(n353) );
  NOR2_X1 U416 ( .A1(n354), .A2(n353), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT46), .B(KEYINPUT105), .Z(n358) );
  XNOR2_X1 U419 ( .A(KEYINPUT41), .B(n572), .ZN(n561) );
  NAND2_X1 U420 ( .A1(n561), .A2(n556), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  NAND2_X1 U422 ( .A1(n359), .A2(n565), .ZN(n360) );
  NOR2_X1 U423 ( .A1(n567), .A2(n360), .ZN(n361) );
  XNOR2_X1 U424 ( .A(KEYINPUT47), .B(n361), .ZN(n362) );
  NAND2_X1 U425 ( .A1(n363), .A2(n362), .ZN(n365) );
  XNOR2_X1 U426 ( .A(KEYINPUT107), .B(KEYINPUT48), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n469) );
  XOR2_X1 U428 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n369) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U431 ( .A(n370), .B(KEYINPUT84), .Z(n372) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n371) );
  XOR2_X1 U433 ( .A(n372), .B(n371), .Z(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U435 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n376) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n422) );
  XNOR2_X1 U438 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n377), .B(G211GAT), .ZN(n417) );
  XNOR2_X1 U440 ( .A(n422), .B(n417), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n516) );
  XNOR2_X1 U442 ( .A(n516), .B(KEYINPUT27), .ZN(n450) );
  XOR2_X1 U443 ( .A(KEYINPUT82), .B(KEYINPUT4), .Z(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT81), .B(KEYINPUT5), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n398) );
  XOR2_X1 U446 ( .A(G85GAT), .B(G148GAT), .Z(n383) );
  XNOR2_X1 U447 ( .A(G29GAT), .B(G162GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U449 ( .A(KEYINPUT6), .B(G57GAT), .Z(n385) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(G155GAT), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U452 ( .A(n387), .B(n386), .Z(n396) );
  XOR2_X1 U453 ( .A(G127GAT), .B(G134GAT), .Z(n389) );
  XNOR2_X1 U454 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(n390), .ZN(n433) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n391), .B(KEYINPUT2), .ZN(n416) );
  XOR2_X1 U459 ( .A(n416), .B(KEYINPUT1), .Z(n393) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U462 ( .A(n433), .B(n394), .Z(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n549) );
  NAND2_X1 U465 ( .A1(n450), .A2(n549), .ZN(n442) );
  NOR2_X1 U466 ( .A1(n469), .A2(n442), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n534) );
  XOR2_X1 U468 ( .A(KEYINPUT79), .B(G78GAT), .Z(n402) );
  NAND2_X1 U469 ( .A1(G228GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U471 ( .A(KEYINPUT24), .B(n403), .ZN(n405) );
  XOR2_X1 U472 ( .A(KEYINPUT22), .B(G218GAT), .Z(n409) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U475 ( .A(KEYINPUT23), .B(G204GAT), .Z(n413) );
  XNOR2_X1 U476 ( .A(KEYINPUT80), .B(KEYINPUT78), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n550) );
  XOR2_X1 U481 ( .A(KEYINPUT75), .B(KEYINPUT20), .Z(n421) );
  XNOR2_X1 U482 ( .A(KEYINPUT77), .B(KEYINPUT76), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n432) );
  XOR2_X1 U484 ( .A(G99GAT), .B(G71GAT), .Z(n424) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U487 ( .A(n425), .B(G190GAT), .Z(n430) );
  XOR2_X1 U488 ( .A(G176GAT), .B(G183GAT), .Z(n427) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n434) );
  INV_X1 U494 ( .A(n554), .ZN(n435) );
  OR2_X1 U495 ( .A1(n520), .A2(n435), .ZN(n436) );
  OR2_X1 U496 ( .A1(n534), .A2(n436), .ZN(n437) );
  INV_X1 U497 ( .A(n529), .ZN(n438) );
  NOR2_X1 U498 ( .A1(n565), .A2(n438), .ZN(n441) );
  NOR2_X1 U499 ( .A1(n520), .A2(n442), .ZN(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT86), .B(n443), .Z(n444) );
  NOR2_X1 U501 ( .A1(n554), .A2(n444), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT87), .ZN(n455) );
  INV_X1 U503 ( .A(n549), .ZN(n466) );
  NAND2_X1 U504 ( .A1(n554), .A2(n516), .ZN(n446) );
  NAND2_X1 U505 ( .A1(n550), .A2(n446), .ZN(n447) );
  XOR2_X1 U506 ( .A(KEYINPUT25), .B(n447), .Z(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT88), .B(KEYINPUT26), .ZN(n449) );
  NOR2_X1 U508 ( .A1(n554), .A2(n550), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n533) );
  NAND2_X1 U510 ( .A1(n533), .A2(n450), .ZN(n451) );
  NAND2_X1 U511 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U512 ( .A1(n466), .A2(n453), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n455), .A2(n454), .ZN(n481) );
  NOR2_X1 U514 ( .A1(n575), .A2(n578), .ZN(n456) );
  AND2_X1 U515 ( .A1(n481), .A2(n456), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n572), .A2(n556), .ZN(n483) );
  NOR2_X1 U517 ( .A1(n513), .A2(n483), .ZN(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT95), .B(KEYINPUT38), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U520 ( .A(KEYINPUT94), .B(n462), .Z(n498) );
  NAND2_X1 U521 ( .A1(n498), .A2(n554), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT40), .B(KEYINPUT97), .Z(n463) );
  NAND2_X1 U523 ( .A1(n466), .A2(n533), .ZN(n472) );
  XNOR2_X1 U524 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT54), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n516), .B(KEYINPUT117), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(n548) );
  OR2_X1 U529 ( .A1(n472), .A2(n548), .ZN(n473) );
  XOR2_X1 U530 ( .A(n473), .B(KEYINPUT124), .Z(n576) );
  NAND2_X1 U531 ( .A1(n576), .A2(n556), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT59), .ZN(n478) );
  XOR2_X1 U535 ( .A(G197GAT), .B(KEYINPUT125), .Z(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(G1352GAT) );
  NOR2_X1 U537 ( .A1(n567), .A2(n479), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n501) );
  NOR2_X1 U540 ( .A1(n483), .A2(n501), .ZN(n491) );
  NAND2_X1 U541 ( .A1(n549), .A2(n491), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  XOR2_X1 U544 ( .A(G8GAT), .B(KEYINPUT89), .Z(n487) );
  NAND2_X1 U545 ( .A1(n491), .A2(n516), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT90), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U548 ( .A1(n491), .A2(n554), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n520), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U553 ( .A1(n498), .A2(n549), .ZN(n494) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT91), .Z(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n496) );
  XOR2_X1 U556 ( .A(KEYINPUT39), .B(KEYINPUT96), .Z(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n498), .A2(n516), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n520), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT98), .B(KEYINPUT42), .Z(n503) );
  NAND2_X1 U563 ( .A1(n500), .A2(n561), .ZN(n512) );
  NOR2_X1 U564 ( .A1(n512), .A2(n501), .ZN(n508) );
  NAND2_X1 U565 ( .A1(n508), .A2(n549), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n504), .Z(G1332GAT) );
  XOR2_X1 U568 ( .A(G64GAT), .B(KEYINPUT99), .Z(n506) );
  NAND2_X1 U569 ( .A1(n508), .A2(n516), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n554), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT100), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n520), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U578 ( .A(KEYINPUT101), .B(n514), .Z(n521) );
  NAND2_X1 U579 ( .A1(n549), .A2(n521), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT102), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n554), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT103), .Z(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n556), .A2(n529), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT110), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n561), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT111), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U597 ( .A1(n529), .A2(n567), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n538) );
  INV_X1 U601 ( .A(n533), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT112), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n546), .A2(n556), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n541) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U610 ( .A(KEYINPUT115), .B(n542), .Z(n544) );
  NAND2_X1 U611 ( .A1(n546), .A2(n561), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U613 ( .A1(n546), .A2(n575), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U615 ( .A1(n546), .A2(n567), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U617 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n564) );
  INV_X1 U622 ( .A(n564), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n568), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(n560), .Z(n563) );
  NAND2_X1 U629 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n571), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n576), .ZN(n579) );
  OR2_X1 U639 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

