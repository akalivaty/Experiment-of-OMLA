

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U548 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  INV_X1 U549 ( .A(KEYINPUT29), .ZN(n708) );
  INV_X1 U550 ( .A(KEYINPUT107), .ZN(n729) );
  XNOR2_X1 U551 ( .A(n735), .B(n734), .ZN(n742) );
  NOR2_X1 U552 ( .A1(G651), .A2(n636), .ZN(n646) );
  NOR2_X2 U553 ( .A1(G2105), .A2(n521), .ZN(n550) );
  NOR2_X1 U554 ( .A1(n766), .A2(n749), .ZN(n514) );
  XNOR2_X1 U555 ( .A(n720), .B(KEYINPUT30), .ZN(n721) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n724) );
  XNOR2_X1 U557 ( .A(n724), .B(KEYINPUT106), .ZN(n725) );
  XNOR2_X1 U558 ( .A(n726), .B(n725), .ZN(n727) );
  INV_X1 U559 ( .A(KEYINPUT32), .ZN(n734) );
  INV_X1 U560 ( .A(n1003), .ZN(n746) );
  NAND2_X1 U561 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U562 ( .A1(G8), .A2(n718), .ZN(n766) );
  NOR2_X1 U563 ( .A1(G543), .A2(n529), .ZN(n530) );
  INV_X1 U564 ( .A(KEYINPUT112), .ZN(n807) );
  XOR2_X1 U565 ( .A(KEYINPUT74), .B(n546), .Z(n993) );
  NOR2_X1 U566 ( .A1(n525), .A2(n524), .ZN(G160) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n515), .Z(n867) );
  NAND2_X1 U568 ( .A1(G137), .A2(n867), .ZN(n516) );
  XNOR2_X1 U569 ( .A(n516), .B(KEYINPUT65), .ZN(n525) );
  INV_X1 U570 ( .A(G2104), .ZN(n521) );
  NAND2_X1 U571 ( .A1(G101), .A2(n550), .ZN(n517) );
  XNOR2_X1 U572 ( .A(n517), .B(KEYINPUT23), .ZN(n520) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U574 ( .A1(G113), .A2(n871), .ZN(n518) );
  XOR2_X1 U575 ( .A(KEYINPUT64), .B(n518), .Z(n519) );
  NOR2_X1 U576 ( .A1(n520), .A2(n519), .ZN(n523) );
  AND2_X1 U577 ( .A1(n521), .A2(G2105), .ZN(n870) );
  NAND2_X1 U578 ( .A1(n870), .A2(G125), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U581 ( .A1(n641), .A2(G90), .ZN(n527) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n636) );
  XOR2_X1 U583 ( .A(KEYINPUT66), .B(G651), .Z(n529) );
  NOR2_X1 U584 ( .A1(n636), .A2(n529), .ZN(n642) );
  NAND2_X1 U585 ( .A1(G77), .A2(n642), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U587 ( .A(KEYINPUT9), .B(n528), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G52), .A2(n646), .ZN(n533) );
  XNOR2_X1 U589 ( .A(n530), .B(KEYINPUT68), .ZN(n531) );
  XOR2_X2 U590 ( .A(KEYINPUT1), .B(n531), .Z(n647) );
  NAND2_X1 U591 ( .A1(G64), .A2(n647), .ZN(n532) );
  AND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n535), .A2(n534), .ZN(G301) );
  INV_X1 U594 ( .A(G301), .ZN(G171) );
  INV_X1 U595 ( .A(G860), .ZN(n591) );
  NAND2_X1 U596 ( .A1(G81), .A2(n641), .ZN(n536) );
  XOR2_X1 U597 ( .A(KEYINPUT12), .B(n536), .Z(n537) );
  XNOR2_X1 U598 ( .A(n537), .B(KEYINPUT73), .ZN(n539) );
  NAND2_X1 U599 ( .A1(G68), .A2(n642), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n540), .B(KEYINPUT13), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G43), .A2(n646), .ZN(n541) );
  AND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n647), .A2(G56), .ZN(n543) );
  XNOR2_X1 U605 ( .A(KEYINPUT14), .B(n543), .ZN(n544) );
  AND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U607 ( .A1(n591), .A2(n993), .ZN(G153) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(n867), .A2(G138), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G126), .A2(n870), .ZN(n547) );
  XOR2_X1 U613 ( .A(KEYINPUT91), .B(n547), .Z(n548) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G102), .A2(n550), .ZN(n552) );
  NAND2_X1 U616 ( .A1(G114), .A2(n871), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n554), .A2(n553), .ZN(G164) );
  NAND2_X1 U619 ( .A1(G51), .A2(n646), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G63), .A2(n647), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(n557), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n641), .A2(G89), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G76), .A2(n642), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(n561), .B(KEYINPUT5), .Z(n562) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT76), .B(n564), .Z(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT7), .B(n565), .ZN(G168) );
  NAND2_X1 U631 ( .A1(G94), .A2(G452), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U635 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n569) );
  INV_X1 U636 ( .A(G223), .ZN(n835) );
  NAND2_X1 U637 ( .A1(G567), .A2(n835), .ZN(n568) );
  XNOR2_X1 U638 ( .A(n569), .B(n568), .ZN(G234) );
  INV_X1 U639 ( .A(G868), .ZN(n661) );
  NOR2_X1 U640 ( .A1(n661), .A2(G171), .ZN(n570) );
  XNOR2_X1 U641 ( .A(n570), .B(KEYINPUT75), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n641), .A2(G92), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G79), .A2(n642), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G54), .A2(n646), .ZN(n574) );
  NAND2_X1 U646 ( .A1(G66), .A2(n647), .ZN(n573) );
  NAND2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U649 ( .A(KEYINPUT15), .B(n577), .Z(n1000) );
  NAND2_X1 U650 ( .A1(n661), .A2(n690), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(G284) );
  XOR2_X1 U652 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U653 ( .A1(G91), .A2(n641), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n580), .B(KEYINPUT70), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n647), .A2(G65), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n646), .A2(G53), .ZN(n584) );
  NAND2_X1 U658 ( .A1(G78), .A2(n642), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n985) );
  XNOR2_X1 U661 ( .A(n985), .B(KEYINPUT71), .ZN(G299) );
  XNOR2_X1 U662 ( .A(KEYINPUT77), .B(G868), .ZN(n587) );
  NOR2_X1 U663 ( .A1(G286), .A2(n587), .ZN(n589) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U666 ( .A(KEYINPUT78), .B(n590), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n592), .A2(n1000), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT79), .ZN(n594) );
  XOR2_X1 U670 ( .A(KEYINPUT16), .B(n594), .Z(G148) );
  NAND2_X1 U671 ( .A1(n1000), .A2(G868), .ZN(n595) );
  NOR2_X1 U672 ( .A1(G559), .A2(n595), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n596), .B(KEYINPUT80), .ZN(n598) );
  NOR2_X1 U674 ( .A1(n993), .A2(G868), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U676 ( .A1(n870), .A2(G123), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n599), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U678 ( .A1(G111), .A2(n871), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G135), .A2(n867), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G99), .A2(n550), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n962) );
  XOR2_X1 U684 ( .A(G2096), .B(n962), .Z(n606) );
  NOR2_X1 U685 ( .A1(G2100), .A2(n606), .ZN(n607) );
  XNOR2_X1 U686 ( .A(KEYINPUT81), .B(n607), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n641), .A2(G93), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G80), .A2(n642), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G55), .A2(n646), .ZN(n611) );
  NAND2_X1 U691 ( .A1(G67), .A2(n647), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n660) );
  NAND2_X1 U694 ( .A1(G559), .A2(n1000), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(n993), .ZN(n658) );
  XNOR2_X1 U696 ( .A(KEYINPUT82), .B(n658), .ZN(n615) );
  NOR2_X1 U697 ( .A1(G860), .A2(n615), .ZN(n616) );
  XOR2_X1 U698 ( .A(n660), .B(n616), .Z(G145) );
  NAND2_X1 U699 ( .A1(n641), .A2(G88), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G75), .A2(n642), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G62), .A2(n647), .ZN(n619) );
  XNOR2_X1 U703 ( .A(KEYINPUT87), .B(n619), .ZN(n620) );
  NOR2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n646), .A2(G50), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(G303) );
  INV_X1 U707 ( .A(G303), .ZN(G166) );
  NAND2_X1 U708 ( .A1(n642), .A2(G73), .ZN(n624) );
  XNOR2_X1 U709 ( .A(n624), .B(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G48), .A2(n646), .ZN(n626) );
  NAND2_X1 U711 ( .A1(G61), .A2(n647), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n641), .A2(G86), .ZN(n627) );
  XOR2_X1 U714 ( .A(KEYINPUT86), .B(n627), .Z(n628) );
  NOR2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U717 ( .A1(n646), .A2(G49), .ZN(n632) );
  XOR2_X1 U718 ( .A(KEYINPUT83), .B(n632), .Z(n634) );
  NAND2_X1 U719 ( .A1(G651), .A2(G74), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U721 ( .A(KEYINPUT84), .B(n635), .Z(n638) );
  NAND2_X1 U722 ( .A1(n636), .A2(G87), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U724 ( .A1(n647), .A2(n639), .ZN(n640) );
  XNOR2_X1 U725 ( .A(KEYINPUT85), .B(n640), .ZN(G288) );
  NAND2_X1 U726 ( .A1(n641), .A2(G85), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G72), .A2(n642), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U729 ( .A(KEYINPUT67), .B(n645), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G47), .A2(n646), .ZN(n649) );
  NAND2_X1 U731 ( .A1(G60), .A2(n647), .ZN(n648) );
  AND2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(G290) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(n660), .ZN(n652) );
  XNOR2_X1 U735 ( .A(G299), .B(n652), .ZN(n653) );
  XNOR2_X1 U736 ( .A(KEYINPUT88), .B(n653), .ZN(n656) );
  XNOR2_X1 U737 ( .A(G166), .B(G305), .ZN(n654) );
  XNOR2_X1 U738 ( .A(n654), .B(G288), .ZN(n655) );
  XNOR2_X1 U739 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U740 ( .A(n657), .B(G290), .ZN(n884) );
  XNOR2_X1 U741 ( .A(n658), .B(n884), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U753 ( .A1(G218), .A2(n669), .ZN(n670) );
  XOR2_X1 U754 ( .A(KEYINPUT89), .B(n670), .Z(n671) );
  NAND2_X1 U755 ( .A1(G96), .A2(n671), .ZN(n840) );
  NAND2_X1 U756 ( .A1(n840), .A2(G2106), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U758 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U759 ( .A1(G108), .A2(n673), .ZN(n839) );
  NAND2_X1 U760 ( .A1(n839), .A2(G567), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n842) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n676) );
  XNOR2_X1 U763 ( .A(KEYINPUT90), .B(n676), .ZN(n677) );
  NOR2_X1 U764 ( .A1(n842), .A2(n677), .ZN(n838) );
  NAND2_X1 U765 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n789) );
  INV_X1 U767 ( .A(n789), .ZN(n678) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n790) );
  NAND2_X2 U769 ( .A1(n678), .A2(n790), .ZN(n718) );
  NOR2_X1 U770 ( .A1(G1971), .A2(n766), .ZN(n680) );
  NOR2_X1 U771 ( .A1(G2090), .A2(n718), .ZN(n679) );
  NOR2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n681), .A2(G303), .ZN(n682) );
  XNOR2_X1 U774 ( .A(KEYINPUT108), .B(n682), .ZN(n732) );
  INV_X1 U775 ( .A(n1000), .ZN(n690) );
  INV_X1 U776 ( .A(n718), .ZN(n683) );
  NAND2_X1 U777 ( .A1(n683), .A2(G1996), .ZN(n684) );
  XNOR2_X1 U778 ( .A(n684), .B(KEYINPUT26), .ZN(n686) );
  NAND2_X1 U779 ( .A1(G1341), .A2(n718), .ZN(n685) );
  NAND2_X1 U780 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n687), .B(KEYINPUT104), .ZN(n688) );
  NOR2_X1 U782 ( .A1(n993), .A2(n688), .ZN(n691) );
  INV_X1 U783 ( .A(n691), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n691), .A2(n1000), .ZN(n695) );
  INV_X1 U786 ( .A(n718), .ZN(n711) );
  NOR2_X1 U787 ( .A1(n711), .A2(G1348), .ZN(n693) );
  NOR2_X1 U788 ( .A1(G2067), .A2(n718), .ZN(n692) );
  NOR2_X1 U789 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n703) );
  NAND2_X1 U792 ( .A1(G1956), .A2(n718), .ZN(n698) );
  XNOR2_X1 U793 ( .A(KEYINPUT103), .B(n698), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n711), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U795 ( .A(KEYINPUT27), .B(n699), .ZN(n700) );
  NOR2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n985), .A2(n704), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n985), .A2(n704), .ZN(n705) );
  XOR2_X1 U800 ( .A(n705), .B(KEYINPUT28), .Z(n706) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U802 ( .A(n709), .B(n708), .ZN(n715) );
  XNOR2_X1 U803 ( .A(KEYINPUT101), .B(G1961), .ZN(n936) );
  NAND2_X1 U804 ( .A1(n718), .A2(n936), .ZN(n710) );
  XNOR2_X1 U805 ( .A(n710), .B(KEYINPUT102), .ZN(n713) );
  XNOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .ZN(n917) );
  NAND2_X1 U807 ( .A1(n711), .A2(n917), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n716), .A2(G171), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n728) );
  OR2_X1 U811 ( .A1(n716), .A2(G171), .ZN(n717) );
  XNOR2_X1 U812 ( .A(n717), .B(KEYINPUT105), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n766), .ZN(n740) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n718), .ZN(n736) );
  NOR2_X1 U815 ( .A1(n740), .A2(n736), .ZN(n719) );
  NAND2_X1 U816 ( .A1(G8), .A2(n719), .ZN(n720) );
  NOR2_X1 U817 ( .A1(G168), .A2(n721), .ZN(n722) );
  NOR2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n738) );
  NAND2_X1 U820 ( .A1(n738), .A2(G286), .ZN(n730) );
  XNOR2_X1 U821 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U823 ( .A1(n733), .A2(G8), .ZN(n735) );
  NAND2_X1 U824 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n759) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n743) );
  XNOR2_X1 U829 ( .A(n743), .B(KEYINPUT109), .ZN(n745) );
  INV_X1 U830 ( .A(KEYINPUT33), .ZN(n744) );
  AND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  OR2_X1 U833 ( .A1(n759), .A2(n748), .ZN(n756) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n988) );
  INV_X1 U835 ( .A(n988), .ZN(n749) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n514), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n750), .A2(n766), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n754) );
  XOR2_X1 U840 ( .A(KEYINPUT110), .B(G1981), .Z(n753) );
  XNOR2_X1 U841 ( .A(G305), .B(n753), .ZN(n990) );
  AND2_X1 U842 ( .A1(n754), .A2(n990), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n763) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n757) );
  XOR2_X1 U845 ( .A(KEYINPUT111), .B(n757), .Z(n758) );
  AND2_X1 U846 ( .A1(G8), .A2(n758), .ZN(n760) );
  OR2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n761), .A2(n766), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n769) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U851 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT100), .ZN(n768) );
  NOR2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n806) );
  NAND2_X1 U855 ( .A1(G129), .A2(n870), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G117), .A2(n871), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U858 ( .A(KEYINPUT96), .B(n772), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G105), .A2(n550), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT38), .ZN(n774) );
  XNOR2_X1 U861 ( .A(n774), .B(KEYINPUT97), .ZN(n775) );
  NOR2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n867), .A2(G141), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n878) );
  NAND2_X1 U865 ( .A1(G1996), .A2(n878), .ZN(n788) );
  XOR2_X1 U866 ( .A(KEYINPUT95), .B(G1991), .Z(n920) );
  NAND2_X1 U867 ( .A1(G131), .A2(n867), .ZN(n779) );
  XNOR2_X1 U868 ( .A(n779), .B(KEYINPUT94), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G119), .A2(n870), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G95), .A2(n550), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G107), .A2(n871), .ZN(n782) );
  XNOR2_X1 U873 ( .A(KEYINPUT93), .B(n782), .ZN(n783) );
  NOR2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n863) );
  NAND2_X1 U876 ( .A1(n920), .A2(n863), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n963) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n820) );
  NAND2_X1 U879 ( .A1(n963), .A2(n820), .ZN(n791) );
  XNOR2_X1 U880 ( .A(n791), .B(KEYINPUT98), .ZN(n809) );
  NAND2_X1 U881 ( .A1(G140), .A2(n867), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G104), .A2(n550), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n794), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G128), .A2(n870), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G116), .A2(n871), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U888 ( .A(KEYINPUT35), .B(n797), .Z(n798) );
  NOR2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U890 ( .A(KEYINPUT36), .B(n800), .Z(n864) );
  XOR2_X1 U891 ( .A(KEYINPUT37), .B(G2067), .Z(n817) );
  AND2_X1 U892 ( .A1(n864), .A2(n817), .ZN(n976) );
  NAND2_X1 U893 ( .A1(n820), .A2(n976), .ZN(n815) );
  NAND2_X1 U894 ( .A1(n809), .A2(n815), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT99), .ZN(n804) );
  XNOR2_X1 U896 ( .A(G1986), .B(KEYINPUT92), .ZN(n802) );
  XNOR2_X1 U897 ( .A(n802), .B(G290), .ZN(n995) );
  NAND2_X1 U898 ( .A1(n995), .A2(n820), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(n807), .ZN(n823) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n878), .ZN(n972) );
  INV_X1 U903 ( .A(n809), .ZN(n812) );
  NOR2_X1 U904 ( .A1(n920), .A2(n863), .ZN(n964) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n964), .A2(n810), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n972), .A2(n813), .ZN(n814) );
  XNOR2_X1 U909 ( .A(KEYINPUT39), .B(n814), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n817), .A2(n864), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT113), .ZN(n981) );
  NAND2_X1 U913 ( .A1(n819), .A2(n981), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n824), .ZN(G329) );
  XNOR2_X1 U917 ( .A(G2454), .B(G2435), .ZN(n833) );
  XNOR2_X1 U918 ( .A(KEYINPUT114), .B(G2427), .ZN(n831) );
  XOR2_X1 U919 ( .A(G2430), .B(G2446), .Z(n826) );
  XNOR2_X1 U920 ( .A(G2443), .B(G2451), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U922 ( .A(n827), .B(G2438), .Z(n829) );
  XNOR2_X1 U923 ( .A(G1348), .B(G1341), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(G14), .ZN(n906) );
  XNOR2_X1 U928 ( .A(KEYINPUT115), .B(n906), .ZN(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U931 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n841), .B(KEYINPUT116), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  INV_X1 U941 ( .A(n842), .ZN(G319) );
  NAND2_X1 U942 ( .A1(G100), .A2(n550), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n843), .B(KEYINPUT118), .ZN(n846) );
  NAND2_X1 U944 ( .A1(G124), .A2(n870), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n844), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U946 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U947 ( .A1(G136), .A2(n867), .ZN(n848) );
  NAND2_X1 U948 ( .A1(G112), .A2(n871), .ZN(n847) );
  NAND2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U950 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U951 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n861) );
  NAND2_X1 U952 ( .A1(G130), .A2(n870), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G118), .A2(n871), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G142), .A2(n867), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G106), .A2(n550), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(KEYINPUT45), .B(n855), .ZN(n856) );
  XNOR2_X1 U959 ( .A(KEYINPUT119), .B(n856), .ZN(n857) );
  NOR2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n962), .B(n859), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n866) );
  XNOR2_X1 U964 ( .A(G160), .B(n864), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n881) );
  NAND2_X1 U966 ( .A1(G139), .A2(n867), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G103), .A2(n550), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G127), .A2(n870), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G115), .A2(n871), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n967) );
  XOR2_X1 U974 ( .A(G162), .B(n967), .Z(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(G164), .B(n879), .Z(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U978 ( .A1(G37), .A2(n882), .ZN(G395) );
  XNOR2_X1 U979 ( .A(G171), .B(n690), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n883), .B(G286), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n993), .B(n884), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U983 ( .A1(G37), .A2(n887), .ZN(G397) );
  XOR2_X1 U984 ( .A(G1956), .B(G1961), .Z(n889) );
  XNOR2_X1 U985 ( .A(G1986), .B(G1966), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U987 ( .A(G1971), .B(G1976), .Z(n891) );
  XNOR2_X1 U988 ( .A(G1996), .B(G1991), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U991 ( .A(KEYINPUT117), .B(G2474), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U993 ( .A(G1981), .B(KEYINPUT41), .Z(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(G229) );
  XOR2_X1 U995 ( .A(G2100), .B(G2096), .Z(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT42), .B(G2678), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U998 ( .A(KEYINPUT43), .B(G2090), .Z(n901) );
  XNOR2_X1 U999 ( .A(G2067), .B(G2072), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G2084), .B(G2078), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(G227) );
  NAND2_X1 U1004 ( .A1(n906), .A2(G319), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(KEYINPUT120), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n908), .B(KEYINPUT121), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n911) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1014 ( .A(G2067), .B(G26), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(G2072), .B(G33), .ZN(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(KEYINPUT124), .B(n916), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G1996), .B(G32), .Z(n919) );
  XNOR2_X1 U1019 ( .A(n917), .B(G27), .ZN(n918) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n924) );
  XOR2_X1 U1021 ( .A(n920), .B(G25), .Z(n921) );
  NAND2_X1 U1022 ( .A1(n921), .A2(G28), .ZN(n922) );
  XOR2_X1 U1023 ( .A(KEYINPUT123), .B(n922), .Z(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n927), .B(KEYINPUT53), .ZN(n930) );
  XOR2_X1 U1027 ( .A(G2084), .B(G34), .Z(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT54), .B(n928), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G35), .B(G2090), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(KEYINPUT125), .B(n933), .Z(n934) );
  NOR2_X1 U1033 ( .A1(G29), .A2(n934), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(n935), .ZN(n1014) );
  XOR2_X1 U1035 ( .A(G16), .B(KEYINPUT126), .Z(n959) );
  XOR2_X1 U1036 ( .A(G1966), .B(G21), .Z(n938) );
  XNOR2_X1 U1037 ( .A(n936), .B(G5), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n956) );
  XNOR2_X1 U1039 ( .A(G1986), .B(G24), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n942) );
  XOR2_X1 U1042 ( .A(G1976), .B(G23), .Z(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(n944), .B(n943), .ZN(n954) );
  XOR2_X1 U1046 ( .A(G1348), .B(KEYINPUT59), .Z(n945) );
  XNOR2_X1 U1047 ( .A(G4), .B(n945), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(G20), .B(G1956), .ZN(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(G1341), .B(G19), .ZN(n948) );
  NOR2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1053 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1054 ( .A(KEYINPUT60), .B(n952), .Z(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(n957), .B(KEYINPUT61), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n960), .ZN(n1012) );
  XOR2_X1 U1060 ( .A(G2084), .B(G160), .Z(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n980) );
  XOR2_X1 U1064 ( .A(G2072), .B(n967), .Z(n969) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n970), .ZN(n978) );
  XOR2_X1 U1068 ( .A(G2090), .B(G162), .Z(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1070 ( .A(KEYINPUT122), .B(n973), .Z(n974) );
  XOR2_X1 U1071 ( .A(KEYINPUT51), .B(n974), .Z(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT52), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n984), .A2(G29), .ZN(n1010) );
  XNOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XOR2_X1 U1079 ( .A(n985), .B(G1956), .Z(n987) );
  XNOR2_X1 U1080 ( .A(G303), .B(G1971), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n999) );
  XNOR2_X1 U1083 ( .A(G168), .B(G1966), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(KEYINPUT57), .B(n992), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n993), .B(G1341), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G171), .B(G1961), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1015), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

