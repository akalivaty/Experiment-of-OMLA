

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n664, n665, n666, n668,
         n669, n670, n671, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779;

  AND2_X1 U379 ( .A1(n358), .A2(n357), .ZN(n664) );
  AND2_X1 U380 ( .A1(n365), .A2(n364), .ZN(n673) );
  AND2_X1 U381 ( .A1(n368), .A2(n367), .ZN(n654) );
  AND2_X1 U382 ( .A1(n371), .A2(n370), .ZN(n688) );
  INV_X1 U383 ( .A(n686), .ZN(n362) );
  INV_X1 U384 ( .A(n686), .ZN(n357) );
  INV_X1 U385 ( .A(n686), .ZN(n364) );
  INV_X1 U386 ( .A(n686), .ZN(n367) );
  INV_X1 U387 ( .A(n686), .ZN(n370) );
  BUF_X1 U388 ( .A(n681), .Z(n390) );
  INV_X1 U389 ( .A(n661), .ZN(n359) );
  AND2_X2 U390 ( .A1(n440), .A2(n411), .ZN(n681) );
  NOR2_X1 U391 ( .A1(n636), .A2(n733), .ZN(n639) );
  AND2_X1 U392 ( .A1(n777), .A2(n621), .ZN(n623) );
  BUF_X1 U393 ( .A(n565), .Z(n373) );
  XNOR2_X1 U394 ( .A(n601), .B(n600), .ZN(n725) );
  AND2_X1 U395 ( .A1(n599), .A2(n598), .ZN(n626) );
  XNOR2_X1 U396 ( .A(n697), .B(n386), .ZN(n565) );
  OR2_X1 U397 ( .A1(n649), .A2(G902), .ZN(n494) );
  XNOR2_X1 U398 ( .A(n512), .B(n511), .ZN(n554) );
  XNOR2_X1 U399 ( .A(n478), .B(n360), .ZN(n480) );
  XNOR2_X1 U400 ( .A(n361), .B(n476), .ZN(n360) );
  XNOR2_X1 U401 ( .A(n419), .B(n508), .ZN(n758) );
  XNOR2_X1 U402 ( .A(n517), .B(n505), .ZN(n419) );
  XNOR2_X1 U403 ( .A(n497), .B(G134), .ZN(n536) );
  BUF_X1 U404 ( .A(G128), .Z(n374) );
  XNOR2_X1 U405 ( .A(G137), .B(KEYINPUT70), .ZN(n763) );
  XNOR2_X1 U406 ( .A(n662), .B(n359), .ZN(n358) );
  INV_X1 U407 ( .A(n477), .ZN(n361) );
  XNOR2_X2 U408 ( .A(n412), .B(n398), .ZN(n635) );
  NOR2_X2 U409 ( .A1(n749), .A2(n393), .ZN(n630) );
  AND2_X1 U410 ( .A1(n363), .A2(n362), .ZN(G66) );
  XNOR2_X1 U411 ( .A(n666), .B(n665), .ZN(n363) );
  XNOR2_X1 U412 ( .A(n671), .B(n366), .ZN(n365) );
  INV_X1 U413 ( .A(n670), .ZN(n366) );
  XNOR2_X1 U414 ( .A(n651), .B(n369), .ZN(n368) );
  INV_X1 U415 ( .A(n650), .ZN(n369) );
  XNOR2_X1 U416 ( .A(n685), .B(n372), .ZN(n371) );
  INV_X1 U417 ( .A(n684), .ZN(n372) );
  XNOR2_X1 U418 ( .A(n486), .B(KEYINPUT73), .ZN(n498) );
  NOR2_X1 U419 ( .A1(G237), .A2(G953), .ZN(n490) );
  NAND2_X1 U420 ( .A1(n394), .A2(n401), .ZN(n644) );
  XNOR2_X1 U421 ( .A(n615), .B(KEYINPUT32), .ZN(n410) );
  XNOR2_X1 U422 ( .A(n463), .B(n462), .ZN(n612) );
  XNOR2_X1 U423 ( .A(n494), .B(G472), .ZN(n562) );
  INV_X1 U424 ( .A(KEYINPUT77), .ZN(n391) );
  OR2_X1 U425 ( .A1(n647), .A2(n644), .ZN(n411) );
  AND2_X1 U426 ( .A1(n377), .A2(n382), .ZN(n381) );
  NAND2_X1 U427 ( .A1(n410), .A2(n657), .ZN(n622) );
  AND2_X1 U428 ( .A1(n582), .A2(n752), .ZN(n425) );
  NOR2_X1 U429 ( .A1(n659), .A2(n779), .ZN(n423) );
  XNOR2_X1 U430 ( .A(n560), .B(KEYINPUT74), .ZN(n561) );
  NAND2_X1 U431 ( .A1(n387), .A2(n692), .ZN(n752) );
  NOR2_X1 U432 ( .A1(n380), .A2(n415), .ZN(n743) );
  XNOR2_X1 U433 ( .A(n388), .B(n570), .ZN(n387) );
  NAND2_X1 U434 ( .A1(n583), .A2(n392), .ZN(n388) );
  NOR2_X1 U435 ( .A1(n572), .A2(n709), .ZN(n515) );
  NAND2_X1 U436 ( .A1(n385), .A2(n626), .ZN(n601) );
  XNOR2_X1 U437 ( .A(n568), .B(KEYINPUT105), .ZN(n583) );
  XNOR2_X1 U438 ( .A(n428), .B(KEYINPUT71), .ZN(n567) );
  INV_X1 U439 ( .A(n565), .ZN(n385) );
  NOR2_X2 U440 ( .A1(n612), .A2(n689), .ZN(n598) );
  INV_X1 U441 ( .A(n612), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n562), .B(KEYINPUT104), .ZN(n616) );
  XNOR2_X1 U443 ( .A(n493), .B(n383), .ZN(n649) );
  XNOR2_X1 U444 ( .A(n384), .B(n492), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n491), .B(n507), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n766), .B(G146), .ZN(n493) );
  NAND2_X1 U447 ( .A1(n509), .A2(n439), .ZN(n400) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n454) );
  XNOR2_X1 U449 ( .A(n450), .B(n449), .ZN(n532) );
  XNOR2_X1 U450 ( .A(n536), .B(n523), .ZN(n766) );
  XNOR2_X1 U451 ( .A(n427), .B(G125), .ZN(n503) );
  AND2_X1 U452 ( .A1(n382), .A2(KEYINPUT65), .ZN(n433) );
  XNOR2_X1 U453 ( .A(n453), .B(KEYINPUT80), .ZN(n379) );
  XNOR2_X1 U454 ( .A(G116), .B(G107), .ZN(n537) );
  XNOR2_X1 U455 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n453) );
  XNOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n378) );
  OR2_X1 U457 ( .A1(n644), .A2(n645), .ZN(n377) );
  NOR2_X1 U458 ( .A1(n644), .A2(n376), .ZN(n438) );
  OR2_X2 U459 ( .A1(n645), .A2(n400), .ZN(n376) );
  NAND2_X1 U460 ( .A1(n377), .A2(n433), .ZN(n432) );
  NOR2_X1 U461 ( .A1(n380), .A2(n724), .ZN(n552) );
  NAND2_X1 U462 ( .A1(n547), .A2(n571), .ZN(n380) );
  INV_X1 U463 ( .A(KEYINPUT2), .ZN(n382) );
  AND2_X1 U464 ( .A1(n373), .A2(n612), .ZN(n613) );
  NAND2_X1 U465 ( .A1(n373), .A2(n375), .ZN(n633) );
  INV_X1 U466 ( .A(n563), .ZN(n386) );
  INV_X1 U467 ( .A(n646), .ZN(n389) );
  XNOR2_X1 U468 ( .A(n431), .B(n447), .ZN(n430) );
  XNOR2_X1 U469 ( .A(n484), .B(n391), .ZN(n395) );
  NAND2_X1 U470 ( .A1(n442), .A2(n441), .ZN(n392) );
  NAND2_X1 U471 ( .A1(n442), .A2(n441), .ZN(n569) );
  XNOR2_X1 U472 ( .A(n569), .B(n556), .ZN(n415) );
  OR2_X1 U473 ( .A1(n629), .A2(n699), .ZN(n445) );
  NOR2_X2 U474 ( .A1(n629), .A2(n610), .ZN(n412) );
  NAND2_X1 U475 ( .A1(n402), .A2(KEYINPUT82), .ZN(n401) );
  XNOR2_X1 U476 ( .A(n503), .B(n426), .ZN(n765) );
  XNOR2_X1 U477 ( .A(G140), .B(KEYINPUT10), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n409) );
  INV_X1 U479 ( .A(KEYINPUT48), .ZN(n420) );
  NAND2_X1 U480 ( .A1(n422), .A2(n424), .ZN(n421) );
  AND2_X1 U481 ( .A1(n561), .A2(n425), .ZN(n424) );
  INV_X1 U482 ( .A(G237), .ZN(n495) );
  XNOR2_X1 U483 ( .A(KEYINPUT3), .B(G119), .ZN(n507) );
  XNOR2_X1 U484 ( .A(n763), .B(G110), .ZN(n476) );
  INV_X1 U485 ( .A(G146), .ZN(n427) );
  INV_X1 U486 ( .A(KEYINPUT33), .ZN(n600) );
  OR2_X2 U487 ( .A1(n415), .A2(n597), .ZN(n413) );
  AND2_X1 U488 ( .A1(n743), .A2(n557), .ZN(n559) );
  XNOR2_X1 U489 ( .A(n423), .B(n446), .ZN(n422) );
  NOR2_X1 U490 ( .A1(KEYINPUT82), .A2(n408), .ZN(n407) );
  INV_X1 U491 ( .A(n656), .ZN(n408) );
  NOR2_X1 U492 ( .A1(n405), .A2(n404), .ZN(n403) );
  INV_X1 U493 ( .A(n655), .ZN(n404) );
  NOR2_X1 U494 ( .A1(n656), .A2(n588), .ZN(n405) );
  XNOR2_X1 U495 ( .A(KEYINPUT5), .B(G137), .ZN(n485) );
  XNOR2_X1 U496 ( .A(G113), .B(G116), .ZN(n487) );
  INV_X1 U497 ( .A(KEYINPUT8), .ZN(n449) );
  NAND2_X1 U498 ( .A1(n769), .A2(G234), .ZN(n450) );
  XNOR2_X1 U499 ( .A(KEYINPUT69), .B(G131), .ZN(n523) );
  NAND2_X1 U500 ( .A1(n612), .A2(n429), .ZN(n428) );
  AND2_X1 U501 ( .A1(n609), .A2(n397), .ZN(n429) );
  NAND2_X1 U502 ( .A1(n616), .A2(n707), .ZN(n431) );
  NOR2_X1 U503 ( .A1(n437), .A2(n399), .ZN(n435) );
  NOR2_X1 U504 ( .A1(n509), .A2(KEYINPUT65), .ZN(n437) );
  NAND2_X1 U505 ( .A1(n439), .A2(KEYINPUT2), .ZN(n436) );
  XOR2_X1 U506 ( .A(G104), .B(G140), .Z(n475) );
  XNOR2_X1 U507 ( .A(KEYINPUT18), .B(KEYINPUT88), .ZN(n496) );
  XNOR2_X1 U508 ( .A(KEYINPUT87), .B(KEYINPUT17), .ZN(n501) );
  NAND2_X1 U509 ( .A1(G237), .A2(G234), .ZN(n471) );
  OR2_X1 U510 ( .A1(n707), .A2(KEYINPUT86), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n531), .B(n530), .ZN(n573) );
  XNOR2_X1 U512 ( .A(n529), .B(n528), .ZN(n530) );
  BUF_X1 U513 ( .A(n554), .Z(n586) );
  BUF_X2 U514 ( .A(n562), .Z(n697) );
  XNOR2_X1 U515 ( .A(KEYINPUT16), .B(G110), .ZN(n506) );
  INV_X1 U516 ( .A(n476), .ZN(n448) );
  NOR2_X1 U517 ( .A1(n769), .A2(G952), .ZN(n686) );
  NOR2_X1 U518 ( .A1(n381), .A2(n414), .ZN(n730) );
  INV_X1 U519 ( .A(KEYINPUT34), .ZN(n602) );
  NOR2_X1 U520 ( .A1(n629), .A2(n628), .ZN(n393) );
  AND2_X1 U521 ( .A1(n406), .A2(n403), .ZN(n394) );
  NAND2_X1 U522 ( .A1(n707), .A2(KEYINPUT86), .ZN(n396) );
  AND2_X1 U523 ( .A1(n473), .A2(n472), .ZN(n397) );
  XOR2_X1 U524 ( .A(n611), .B(KEYINPUT22), .Z(n398) );
  AND2_X1 U525 ( .A1(n509), .A2(n436), .ZN(n399) );
  INV_X1 U526 ( .A(KEYINPUT82), .ZN(n588) );
  NOR2_X2 U527 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U528 ( .A(n409), .ZN(n402) );
  NAND2_X1 U529 ( .A1(n409), .A2(n407), .ZN(n406) );
  XNOR2_X1 U530 ( .A(n410), .B(G119), .ZN(G21) );
  INV_X1 U531 ( .A(n411), .ZN(n414) );
  XNOR2_X2 U532 ( .A(n413), .B(KEYINPUT0), .ZN(n629) );
  OR2_X2 U533 ( .A1(n683), .A2(n509), .ZN(n512) );
  XNOR2_X1 U534 ( .A(n416), .B(n758), .ZN(n683) );
  XNOR2_X1 U535 ( .A(n417), .B(n418), .ZN(n416) );
  XNOR2_X1 U536 ( .A(n498), .B(n503), .ZN(n417) );
  XNOR2_X1 U537 ( .A(n502), .B(n499), .ZN(n418) );
  NAND2_X1 U538 ( .A1(n434), .A2(n432), .ZN(n440) );
  XNOR2_X2 U539 ( .A(G143), .B(G128), .ZN(n497) );
  NAND2_X1 U540 ( .A1(n395), .A2(n430), .ZN(n572) );
  NOR2_X1 U541 ( .A1(n438), .A2(n435), .ZN(n434) );
  INV_X1 U542 ( .A(KEYINPUT65), .ZN(n439) );
  OR2_X1 U543 ( .A1(n554), .A2(n396), .ZN(n441) );
  AND2_X2 U544 ( .A1(n444), .A2(n443), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n554), .A2(n555), .ZN(n444) );
  XNOR2_X2 U546 ( .A(n445), .B(KEYINPUT31), .ZN(n749) );
  NAND2_X1 U547 ( .A1(n681), .A2(G478), .ZN(n662) );
  XOR2_X1 U548 ( .A(n553), .B(KEYINPUT64), .Z(n446) );
  XOR2_X1 U549 ( .A(KEYINPUT106), .B(KEYINPUT30), .Z(n447) );
  XNOR2_X1 U550 ( .A(n765), .B(n448), .ZN(n457) );
  INV_X1 U551 ( .A(n660), .ZN(n661) );
  XNOR2_X1 U552 ( .A(KEYINPUT36), .B(KEYINPUT109), .ZN(n570) );
  INV_X1 U553 ( .A(KEYINPUT63), .ZN(n653) );
  INV_X4 U554 ( .A(G953), .ZN(n769) );
  NAND2_X1 U555 ( .A1(G221), .A2(n532), .ZN(n452) );
  XNOR2_X1 U556 ( .A(n374), .B(G119), .ZN(n451) );
  XNOR2_X1 U557 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U558 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U559 ( .A(n457), .B(n456), .ZN(n665) );
  INV_X1 U560 ( .A(G902), .ZN(n541) );
  NAND2_X1 U561 ( .A1(n665), .A2(n541), .ZN(n463) );
  XNOR2_X1 U562 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  NAND2_X1 U563 ( .A1(G234), .A2(n643), .ZN(n458) );
  XNOR2_X1 U564 ( .A(KEYINPUT20), .B(n458), .ZN(n464) );
  NAND2_X1 U565 ( .A1(G217), .A2(n464), .ZN(n461) );
  INV_X1 U566 ( .A(KEYINPUT79), .ZN(n459) );
  XNOR2_X1 U567 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U569 ( .A1(n464), .A2(G221), .ZN(n468) );
  XOR2_X1 U570 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n466) );
  INV_X1 U571 ( .A(KEYINPUT93), .ZN(n465) );
  XNOR2_X1 U572 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n468), .B(n467), .ZN(n609) );
  INV_X1 U574 ( .A(n609), .ZN(n689) );
  NOR2_X1 U575 ( .A1(G900), .A2(n769), .ZN(n469) );
  NAND2_X1 U576 ( .A1(n469), .A2(G902), .ZN(n470) );
  NAND2_X1 U577 ( .A1(G952), .A2(n769), .ZN(n594) );
  NAND2_X1 U578 ( .A1(n470), .A2(n594), .ZN(n473) );
  XOR2_X1 U579 ( .A(n471), .B(KEYINPUT14), .Z(n720) );
  INV_X1 U580 ( .A(n720), .ZN(n472) );
  NAND2_X1 U581 ( .A1(G227), .A2(n769), .ZN(n474) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X2 U583 ( .A(KEYINPUT4), .B(G101), .ZN(n486) );
  XNOR2_X1 U584 ( .A(n498), .B(G107), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n493), .B(n480), .ZN(n677) );
  NAND2_X1 U586 ( .A1(n677), .A2(n541), .ZN(n482) );
  XNOR2_X1 U587 ( .A(KEYINPUT72), .B(G469), .ZN(n481) );
  XNOR2_X2 U588 ( .A(n482), .B(n481), .ZN(n571) );
  AND2_X1 U589 ( .A1(n397), .A2(n571), .ZN(n483) );
  AND2_X1 U590 ( .A1(n598), .A2(n483), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n486), .B(n485), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n487), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U593 ( .A(n489), .B(n488), .ZN(n492) );
  XNOR2_X1 U594 ( .A(KEYINPUT76), .B(n490), .ZN(n519) );
  NAND2_X1 U595 ( .A1(n519), .A2(G210), .ZN(n491) );
  NAND2_X1 U596 ( .A1(n541), .A2(n495), .ZN(n510) );
  NAND2_X1 U597 ( .A1(n510), .A2(G214), .ZN(n707) );
  XNOR2_X1 U598 ( .A(n497), .B(n496), .ZN(n499) );
  NAND2_X1 U599 ( .A1(n769), .A2(G224), .ZN(n500) );
  XNOR2_X1 U600 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X2 U601 ( .A(G122), .B(G113), .ZN(n504) );
  XNOR2_X2 U602 ( .A(n504), .B(G104), .ZN(n517) );
  INV_X1 U603 ( .A(n537), .ZN(n505) );
  XNOR2_X1 U604 ( .A(n507), .B(n506), .ZN(n508) );
  INV_X1 U605 ( .A(n643), .ZN(n509) );
  NAND2_X1 U606 ( .A1(n510), .A2(G210), .ZN(n511) );
  XNOR2_X1 U607 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n586), .B(n513), .ZN(n709) );
  XNOR2_X1 U609 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n514) );
  XNOR2_X1 U610 ( .A(n515), .B(n514), .ZN(n589) );
  XOR2_X1 U611 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n516) );
  XNOR2_X1 U612 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n765), .B(n518), .ZN(n527) );
  NAND2_X1 U614 ( .A1(n519), .A2(G214), .ZN(n521) );
  XNOR2_X1 U615 ( .A(KEYINPUT97), .B(KEYINPUT11), .ZN(n520) );
  XNOR2_X1 U616 ( .A(n521), .B(n520), .ZN(n525) );
  XNOR2_X1 U617 ( .A(G143), .B(KEYINPUT99), .ZN(n522) );
  XNOR2_X1 U618 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U619 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n527), .B(n526), .ZN(n669) );
  NOR2_X1 U621 ( .A1(G902), .A2(n669), .ZN(n531) );
  XNOR2_X1 U622 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n529) );
  INV_X1 U623 ( .A(G475), .ZN(n528) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n534) );
  NAND2_X1 U625 ( .A1(G217), .A2(n532), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U627 ( .A(n535), .B(KEYINPUT7), .Z(n540) );
  XNOR2_X1 U628 ( .A(n537), .B(G122), .ZN(n538) );
  XNOR2_X1 U629 ( .A(n536), .B(n538), .ZN(n539) );
  XNOR2_X1 U630 ( .A(n540), .B(n539), .ZN(n660) );
  AND2_X1 U631 ( .A1(n660), .A2(n541), .ZN(n543) );
  XOR2_X1 U632 ( .A(G478), .B(KEYINPUT102), .Z(n542) );
  XNOR2_X1 U633 ( .A(n543), .B(n542), .ZN(n574) );
  OR2_X1 U634 ( .A1(n573), .A2(n574), .ZN(n564) );
  NOR2_X1 U635 ( .A1(n589), .A2(n564), .ZN(n544) );
  XNOR2_X1 U636 ( .A(n544), .B(KEYINPUT40), .ZN(n659) );
  NAND2_X1 U637 ( .A1(n567), .A2(n616), .ZN(n546) );
  INV_X1 U638 ( .A(KEYINPUT28), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n546), .B(n545), .ZN(n547) );
  INV_X1 U640 ( .A(n574), .ZN(n548) );
  AND2_X1 U641 ( .A1(n573), .A2(n548), .ZN(n706) );
  NAND2_X1 U642 ( .A1(n706), .A2(n707), .ZN(n549) );
  NOR2_X1 U643 ( .A1(n549), .A2(n709), .ZN(n551) );
  XNOR2_X1 U644 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n550) );
  XNOR2_X1 U645 ( .A(n551), .B(n550), .ZN(n724) );
  XNOR2_X1 U646 ( .A(n552), .B(KEYINPUT42), .ZN(n779) );
  XNOR2_X1 U647 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n553) );
  INV_X1 U648 ( .A(KEYINPUT86), .ZN(n555) );
  XNOR2_X1 U649 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n556) );
  XOR2_X1 U650 ( .A(KEYINPUT68), .B(KEYINPUT47), .Z(n557) );
  INV_X1 U651 ( .A(n564), .ZN(n745) );
  AND2_X1 U652 ( .A1(n573), .A2(n574), .ZN(n748) );
  NOR2_X1 U653 ( .A1(n745), .A2(n748), .ZN(n579) );
  XOR2_X1 U654 ( .A(n579), .B(KEYINPUT81), .Z(n631) );
  INV_X1 U655 ( .A(n631), .ZN(n558) );
  NAND2_X1 U656 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U657 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n563) );
  NOR2_X1 U658 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U659 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U660 ( .A(n571), .B(KEYINPUT1), .ZN(n599) );
  BUF_X1 U661 ( .A(n599), .Z(n692) );
  INV_X1 U662 ( .A(n572), .ZN(n577) );
  INV_X1 U663 ( .A(n573), .ZN(n575) );
  NAND2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n604) );
  NOR2_X1 U665 ( .A1(n604), .A2(n586), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U667 ( .A(KEYINPUT107), .B(n578), .Z(n778) );
  INV_X1 U668 ( .A(n579), .ZN(n708) );
  NAND2_X1 U669 ( .A1(n743), .A2(n708), .ZN(n580) );
  NAND2_X1 U670 ( .A1(n580), .A2(KEYINPUT47), .ZN(n581) );
  AND2_X1 U671 ( .A1(n778), .A2(n581), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n583), .A2(n707), .ZN(n584) );
  NOR2_X1 U673 ( .A1(n692), .A2(n584), .ZN(n585) );
  XOR2_X1 U674 ( .A(KEYINPUT43), .B(n585), .Z(n587) );
  NAND2_X1 U675 ( .A1(n587), .A2(n586), .ZN(n656) );
  INV_X1 U676 ( .A(n589), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n590), .A2(n748), .ZN(n655) );
  NOR2_X1 U678 ( .A1(G898), .A2(n769), .ZN(n591) );
  XOR2_X1 U679 ( .A(KEYINPUT89), .B(n591), .Z(n759) );
  NAND2_X1 U680 ( .A1(G902), .A2(n759), .ZN(n592) );
  NOR2_X1 U681 ( .A1(n720), .A2(n592), .ZN(n593) );
  XNOR2_X1 U682 ( .A(n593), .B(KEYINPUT90), .ZN(n596) );
  NOR2_X1 U683 ( .A1(n720), .A2(n594), .ZN(n595) );
  NOR2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U685 ( .A1(n629), .A2(n725), .ZN(n603) );
  XNOR2_X1 U686 ( .A(n603), .B(n602), .ZN(n605) );
  XNOR2_X2 U687 ( .A(n606), .B(KEYINPUT35), .ZN(n777) );
  NAND2_X1 U688 ( .A1(n777), .A2(KEYINPUT85), .ZN(n608) );
  INV_X1 U689 ( .A(KEYINPUT44), .ZN(n607) );
  NAND2_X1 U690 ( .A1(n608), .A2(n607), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n706), .A2(n609), .ZN(n610) );
  INV_X1 U692 ( .A(KEYINPUT66), .ZN(n611) );
  AND2_X1 U693 ( .A1(n613), .A2(n692), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n635), .A2(n614), .ZN(n615) );
  OR2_X1 U695 ( .A1(n616), .A2(n375), .ZN(n617) );
  NOR2_X1 U696 ( .A1(n692), .A2(n617), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n635), .A2(n618), .ZN(n657) );
  INV_X1 U698 ( .A(n622), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n625) );
  NOR2_X1 U700 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n641) );
  NAND2_X1 U703 ( .A1(n626), .A2(n697), .ZN(n699) );
  NAND2_X1 U704 ( .A1(n571), .A2(n598), .ZN(n627) );
  OR2_X1 U705 ( .A1(n627), .A2(n697), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n630), .B(KEYINPUT96), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n636) );
  NOR2_X1 U708 ( .A1(n692), .A2(n633), .ZN(n634) );
  AND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n733) );
  INV_X1 U710 ( .A(n777), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n637), .A2(KEYINPUT44), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(KEYINPUT45), .ZN(n645) );
  INV_X1 U715 ( .A(n645), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n646), .A2(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n681), .A2(G472), .ZN(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n654), .B(n653), .ZN(G57) );
  XNOR2_X1 U721 ( .A(n655), .B(G134), .ZN(G36) );
  XNOR2_X1 U722 ( .A(n656), .B(G140), .ZN(G42) );
  XNOR2_X1 U723 ( .A(n657), .B(G110), .ZN(G12) );
  XNOR2_X1 U724 ( .A(G131), .B(KEYINPUT127), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n659), .B(n658), .ZN(G33) );
  XNOR2_X1 U726 ( .A(n664), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U727 ( .A1(n390), .A2(G217), .ZN(n666) );
  NAND2_X1 U728 ( .A1(n681), .A2(G475), .ZN(n671) );
  XNOR2_X1 U729 ( .A(KEYINPUT67), .B(KEYINPUT59), .ZN(n668) );
  XNOR2_X1 U730 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U731 ( .A(n673), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U732 ( .A1(n390), .A2(G469), .ZN(n679) );
  XOR2_X1 U733 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n675) );
  XNOR2_X1 U734 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U736 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U737 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U738 ( .A1(n680), .A2(n686), .ZN(G54) );
  NAND2_X1 U739 ( .A1(n681), .A2(G210), .ZN(n685) );
  XOR2_X1 U740 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(n688), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U743 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n719) );
  NAND2_X1 U744 ( .A1(n689), .A2(n612), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(KEYINPUT115), .ZN(n691) );
  XNOR2_X1 U746 ( .A(KEYINPUT49), .B(n691), .ZN(n696) );
  NOR2_X1 U747 ( .A1(n598), .A2(n692), .ZN(n693) );
  XOR2_X1 U748 ( .A(KEYINPUT116), .B(n693), .Z(n694) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n694), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n696), .A2(n695), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n698), .A2(n697), .ZN(n701) );
  INV_X1 U752 ( .A(n699), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U754 ( .A(KEYINPUT51), .B(n702), .Z(n703) );
  NOR2_X1 U755 ( .A1(n724), .A2(n703), .ZN(n716) );
  INV_X1 U756 ( .A(n707), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n709), .A2(n704), .ZN(n705) );
  AND2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n713) );
  NAND2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U761 ( .A(KEYINPUT117), .B(n711), .Z(n712) );
  NOR2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n714), .A2(n725), .ZN(n715) );
  NOR2_X1 U764 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U765 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  XNOR2_X1 U766 ( .A(n719), .B(n718), .ZN(n721) );
  NOR2_X1 U767 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U768 ( .A1(n722), .A2(G952), .ZN(n723) );
  XNOR2_X1 U769 ( .A(n723), .B(KEYINPUT120), .ZN(n728) );
  NOR2_X1 U770 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U771 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U772 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U773 ( .A1(n730), .A2(n729), .ZN(n732) );
  XOR2_X1 U774 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n731) );
  XNOR2_X1 U775 ( .A(n732), .B(n731), .ZN(G75) );
  XOR2_X1 U776 ( .A(G101), .B(n733), .Z(G3) );
  NAND2_X1 U777 ( .A1(n393), .A2(n745), .ZN(n734) );
  XNOR2_X1 U778 ( .A(n734), .B(G104), .ZN(G6) );
  XOR2_X1 U779 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n736) );
  NAND2_X1 U780 ( .A1(n393), .A2(n748), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n736), .B(n735), .ZN(n738) );
  XOR2_X1 U782 ( .A(G107), .B(KEYINPUT111), .Z(n737) );
  XNOR2_X1 U783 ( .A(n738), .B(n737), .ZN(G9) );
  XOR2_X1 U784 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n740) );
  NAND2_X1 U785 ( .A1(n743), .A2(n748), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n740), .B(n739), .ZN(n742) );
  XOR2_X1 U787 ( .A(n374), .B(KEYINPUT112), .Z(n741) );
  XNOR2_X1 U788 ( .A(n742), .B(n741), .ZN(G30) );
  NAND2_X1 U789 ( .A1(n743), .A2(n745), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(G146), .ZN(G48) );
  NAND2_X1 U791 ( .A1(n749), .A2(n745), .ZN(n746) );
  XNOR2_X1 U792 ( .A(n746), .B(KEYINPUT114), .ZN(n747) );
  XNOR2_X1 U793 ( .A(G113), .B(n747), .ZN(G15) );
  NAND2_X1 U794 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U795 ( .A(n750), .B(G116), .ZN(G18) );
  XOR2_X1 U796 ( .A(G125), .B(KEYINPUT37), .Z(n751) );
  XNOR2_X1 U797 ( .A(n752), .B(n751), .ZN(G27) );
  NOR2_X1 U798 ( .A1(n389), .A2(G953), .ZN(n757) );
  NAND2_X1 U799 ( .A1(G953), .A2(G224), .ZN(n753) );
  XNOR2_X1 U800 ( .A(KEYINPUT61), .B(n753), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n754), .A2(G898), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n755), .B(KEYINPUT125), .ZN(n756) );
  NOR2_X1 U803 ( .A1(n757), .A2(n756), .ZN(n762) );
  XOR2_X1 U804 ( .A(G101), .B(n758), .Z(n760) );
  NOR2_X1 U805 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U806 ( .A(n762), .B(n761), .Z(G69) );
  XNOR2_X1 U807 ( .A(n763), .B(KEYINPUT4), .ZN(n764) );
  XNOR2_X1 U808 ( .A(n765), .B(n764), .ZN(n768) );
  INV_X1 U809 ( .A(n766), .ZN(n767) );
  XNOR2_X1 U810 ( .A(n768), .B(n767), .ZN(n772) );
  XNOR2_X1 U811 ( .A(n644), .B(n772), .ZN(n770) );
  NAND2_X1 U812 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U813 ( .A(n771), .B(KEYINPUT126), .ZN(n776) );
  XNOR2_X1 U814 ( .A(G227), .B(n772), .ZN(n773) );
  NAND2_X1 U815 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U816 ( .A1(G953), .A2(n774), .ZN(n775) );
  NAND2_X1 U817 ( .A1(n776), .A2(n775), .ZN(G72) );
  XNOR2_X1 U818 ( .A(n777), .B(G122), .ZN(G24) );
  XNOR2_X1 U819 ( .A(G143), .B(n778), .ZN(G45) );
  XOR2_X1 U820 ( .A(G137), .B(n779), .Z(G39) );
endmodule

