//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n207), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n218), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n230), .B(new_n231), .Z(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n223), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n245), .A2(new_n247), .B1(G150), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n249), .A2(KEYINPUT66), .B1(new_n203), .B2(G20), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(KEYINPUT66), .B2(new_n249), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n222), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n253), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n209), .B1(new_n255), .B2(G20), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(new_n259), .B1(new_n209), .B2(new_n257), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT9), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G274), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  INV_X1    g0075(.A(G77), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1698), .B1(new_n271), .B2(new_n272), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(G222), .B2(new_n278), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n268), .B1(new_n210), .B2(new_n270), .C1(new_n279), .C2(new_n265), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(G200), .B2(new_n280), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n262), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT10), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT10), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n262), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n248), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n289), .A2(new_n209), .B1(new_n223), .B2(G68), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n246), .A2(new_n276), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n253), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT11), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n256), .A2(G68), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT12), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n297), .B(new_n298), .C1(new_n295), .C2(new_n294), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n258), .B(G68), .C1(G1), .C2(new_n223), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT14), .ZN(new_n302));
  INV_X1    g0102(.A(G238), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n268), .B1(new_n270), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n229), .A2(G1698), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(G226), .B2(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n305), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n265), .B1(new_n309), .B2(new_n310), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT13), .B1(new_n316), .B2(new_n304), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n302), .B1(new_n318), .B2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT14), .B(new_n320), .C1(new_n315), .C2(new_n317), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(G179), .A3(new_n317), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n315), .A2(KEYINPUT70), .A3(new_n317), .A4(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n322), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(new_n322), .B2(new_n328), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n301), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(new_n247), .B1(G20), .B2(G77), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n244), .B(KEYINPUT67), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n289), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n253), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n276), .B1(new_n255), .B2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n258), .A2(new_n339), .B1(new_n276), .B2(new_n257), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n312), .A2(new_n267), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G244), .ZN(new_n343));
  INV_X1    g0143(.A(G107), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n274), .A2(new_n303), .B1(new_n344), .B2(new_n273), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G232), .B2(new_n278), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n268), .B(new_n343), .C1(new_n346), .C2(new_n265), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n320), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n320), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n338), .A2(new_n340), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n347), .A2(G179), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n349), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n280), .A2(new_n320), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n261), .C1(G179), .C2(new_n280), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n341), .B1(new_n281), .B2(new_n347), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n347), .A2(G200), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n357), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n318), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G190), .ZN(new_n367));
  INV_X1    g0167(.A(new_n301), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n366), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n288), .A2(new_n332), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  INV_X1    g0172(.A(G68), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n202), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n248), .A2(G159), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n271), .A2(new_n223), .A3(new_n272), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n272), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n381), .B1(new_n386), .B2(G68), .ZN(new_n387));
  AOI211_X1 g0187(.A(KEYINPUT72), .B(new_n373), .C1(new_n384), .C2(new_n385), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT16), .B(new_n380), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  XOR2_X1   g0189(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n390));
  NAND2_X1  g0190(.A1(new_n375), .A2(new_n377), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n373), .B1(new_n384), .B2(new_n385), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(new_n396), .A3(new_n253), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n244), .B1(new_n255), .B2(G20), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n258), .B1(new_n257), .B2(new_n244), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n268), .B1(new_n270), .B2(new_n229), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n210), .A2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G223), .B2(G1698), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n307), .A2(new_n308), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n403), .A2(new_n404), .B1(new_n263), .B2(new_n211), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n405), .B2(new_n312), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n406), .A2(new_n320), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n400), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G200), .B2(new_n406), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n397), .A2(new_n399), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT17), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n400), .A2(new_n419), .A3(new_n409), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n397), .A2(new_n399), .A3(new_n416), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n411), .A2(new_n418), .A3(new_n420), .A4(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n371), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G1698), .ZN(new_n426));
  OAI211_X1 g0226(.A(G244), .B(new_n426), .C1(new_n307), .C2(new_n308), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G283), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n429), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n312), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT5), .B(G41), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n266), .A2(G1), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(G257), .A3(new_n265), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(new_n265), .A3(G274), .A4(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n312), .B2(new_n433), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT76), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(G200), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n256), .A2(G97), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n255), .A2(G33), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n222), .A2(new_n256), .A3(new_n252), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(G97), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT7), .B1(new_n404), .B2(new_n223), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n307), .A2(new_n308), .A3(new_n383), .A4(G20), .ZN(new_n454));
  OAI21_X1  g0254(.A(G107), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n289), .A2(new_n276), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT6), .ZN(new_n457));
  AND2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  NOR2_X1   g0258(.A1(G97), .A2(G107), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n344), .A2(KEYINPUT6), .A3(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n456), .B1(new_n462), .B2(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n452), .B1(new_n464), .B2(new_n253), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n434), .A2(G190), .A3(new_n441), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT77), .ZN(new_n469));
  INV_X1    g0269(.A(new_n253), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n455), .B2(new_n463), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n452), .ZN(new_n472));
  INV_X1    g0272(.A(new_n456), .ZN(new_n473));
  XNOR2_X1  g0273(.A(G97), .B(G107), .ZN(new_n474));
  INV_X1    g0274(.A(G97), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n457), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n474), .A2(new_n457), .B1(new_n344), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n477), .B2(new_n223), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n344), .B1(new_n384), .B2(new_n385), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n253), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(KEYINPUT77), .A3(new_n451), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n434), .A2(G179), .A3(new_n441), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n320), .B2(new_n445), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n447), .A2(new_n468), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n303), .A2(G1698), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n307), .B2(new_n308), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT78), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n263), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT78), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n486), .B(new_n493), .C1(new_n308), .C2(new_n307), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n488), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n312), .ZN(new_n496));
  INV_X1    g0296(.A(G179), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n436), .A2(new_n212), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n265), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n265), .A2(G274), .ZN(new_n500));
  INV_X1    g0300(.A(new_n436), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n503), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n223), .B1(new_n310), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n459), .A2(new_n211), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n223), .B(G68), .C1(new_n307), .C2(new_n308), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n506), .B1(new_n246), .B2(new_n475), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(new_n253), .B1(new_n257), .B2(new_n333), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n450), .A2(new_n334), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n505), .A2(new_n320), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n450), .A2(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n505), .B2(G200), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n496), .A2(G190), .A3(new_n503), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n504), .A2(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n485), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n273), .A2(G264), .A3(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(new_n426), .C1(new_n307), .C2(new_n308), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n404), .A2(G303), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n312), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n312), .B1(new_n436), .B2(new_n435), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n435), .A2(new_n436), .ZN(new_n528));
  INV_X1    g0328(.A(G274), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n312), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n527), .A2(G270), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n450), .A2(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n257), .A2(new_n489), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n252), .A2(new_n222), .B1(G20), .B2(new_n489), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n431), .B(new_n223), .C1(G33), .C2(new_n475), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n535), .A2(KEYINPUT20), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT20), .B1(new_n535), .B2(new_n536), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n533), .B(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n532), .A2(KEYINPUT21), .A3(G169), .A4(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(G179), .A3(new_n526), .A4(new_n531), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n532), .A2(G169), .A3(new_n539), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n532), .A2(G200), .ZN(new_n546));
  INV_X1    g0346(.A(new_n539), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(new_n414), .C2(new_n532), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n542), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n223), .B(G87), .C1(new_n307), .C2(new_n308), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT22), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n552), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n273), .A2(new_n554), .A3(new_n223), .A4(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n223), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n344), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n560), .B1(new_n490), .B2(new_n223), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n557), .B1(new_n556), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n253), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n256), .B2(G107), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n256), .A2(new_n565), .A3(G107), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n566), .A2(new_n568), .B1(new_n450), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n437), .A2(G264), .A3(new_n265), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT80), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n527), .A2(KEYINPUT80), .A3(G264), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n273), .A2(G250), .A3(new_n426), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n572), .A2(new_n573), .B1(new_n577), .B2(new_n312), .ZN(new_n578));
  AOI21_X1  g0378(.A(G200), .B1(new_n578), .B2(new_n439), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n577), .A2(new_n312), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n570), .A2(new_n439), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n580), .A2(new_n581), .A3(G190), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n564), .B(new_n569), .C1(new_n579), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n564), .A2(new_n569), .ZN(new_n584));
  OAI21_X1  g0384(.A(G169), .B1(new_n580), .B2(new_n581), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n572), .A2(new_n573), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n577), .A2(new_n312), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(G179), .A3(new_n439), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n521), .A2(new_n549), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n425), .A2(new_n592), .ZN(G372));
  INV_X1    g0393(.A(new_n359), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT81), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n288), .B(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n370), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n357), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n328), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n314), .B1(new_n305), .B2(new_n313), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n316), .A2(new_n304), .A3(KEYINPUT13), .ZN(new_n601));
  OAI21_X1  g0401(.A(G169), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT14), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n318), .A2(new_n302), .A3(G169), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT71), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n368), .B1(new_n606), .B2(new_n329), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n423), .B(new_n418), .C1(new_n598), .C2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n411), .A3(new_n420), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n594), .B1(new_n596), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n583), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n545), .A2(new_n541), .A3(new_n540), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n564), .A2(new_n569), .B1(new_n585), .B2(new_n588), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n521), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n442), .A2(G169), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n465), .B1(new_n617), .B2(new_n483), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n520), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n512), .A2(new_n253), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n333), .A2(new_n257), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n514), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n502), .B1(new_n495), .B2(new_n312), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n504), .B(new_n622), .C1(G169), .C2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n620), .A2(new_n621), .A3(new_n516), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n519), .B(new_n625), .C1(new_n369), .C2(new_n623), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n482), .A2(new_n624), .A3(new_n626), .A4(new_n484), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n619), .A2(new_n628), .A3(new_n624), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n615), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n425), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n610), .A2(new_n631), .ZN(G369));
  NAND3_X1  g0432(.A1(new_n255), .A2(new_n223), .A3(G13), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT82), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(new_n547), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n612), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n549), .B2(new_n639), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n638), .B1(new_n564), .B2(new_n569), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n591), .A2(new_n643), .B1(new_n590), .B2(new_n638), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n591), .ZN(new_n646));
  INV_X1    g0446(.A(new_n638), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n542), .B2(new_n545), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n646), .A2(new_n648), .B1(new_n613), .B2(new_n638), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n649), .ZN(G399));
  NAND2_X1  g0450(.A1(new_n219), .A2(new_n264), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G1), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n508), .A2(G116), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT83), .Z(new_n654));
  OAI22_X1  g0454(.A1(new_n652), .A2(new_n654), .B1(new_n225), .B2(new_n651), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT85), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n624), .B1(new_n627), .B2(KEYINPUT26), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n616), .B1(new_n520), .B2(new_n618), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n369), .B1(new_n442), .B2(new_n443), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n467), .B1(new_n446), .B2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n617), .A2(new_n483), .B1(new_n472), .B2(new_n481), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n625), .B1(new_n623), .B2(new_n369), .ZN(new_n665));
  INV_X1    g0465(.A(new_n519), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n622), .B1(new_n623), .B2(G169), .ZN(new_n667));
  AOI211_X1 g0467(.A(G179), .B(new_n502), .C1(new_n495), .C2(new_n312), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n663), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT86), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n612), .B2(new_n613), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n590), .A2(new_n542), .A3(KEYINPUT86), .A4(new_n545), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n670), .A2(new_n583), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n520), .A2(new_n616), .A3(new_n664), .ZN(new_n675));
  INV_X1    g0475(.A(new_n465), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n484), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT26), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n675), .A2(new_n678), .A3(KEYINPUT85), .A4(new_n624), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n661), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n657), .B1(new_n680), .B2(new_n638), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n657), .B(new_n638), .C1(new_n615), .C2(new_n629), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n532), .A2(new_n497), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n445), .A3(new_n623), .A4(new_n578), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT84), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n578), .A2(new_n439), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n505), .A2(new_n497), .A3(new_n532), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n692), .A2(new_n693), .A3(new_n445), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n690), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n685), .B1(new_n695), .B2(new_n638), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n687), .A2(new_n688), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n697), .B2(KEYINPUT30), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n591), .A2(new_n549), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n670), .A3(new_n638), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n696), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n684), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n656), .B1(new_n707), .B2(G1), .ZN(G364));
  INV_X1    g0508(.A(new_n641), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n641), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT87), .ZN(new_n713));
  INV_X1    g0513(.A(new_n651), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n223), .A2(G13), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n255), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n651), .A2(KEYINPUT87), .A3(new_n716), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n711), .A2(new_n712), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n720), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n207), .A2(G13), .A3(new_n404), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G355), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G116), .B2(new_n219), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n219), .A2(new_n404), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n266), .B2(new_n226), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n239), .A2(G45), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT88), .Z(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n222), .B1(G20), .B2(new_n320), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n722), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n497), .A2(new_n369), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT91), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n223), .A3(G190), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT32), .Z(new_n741));
  INV_X1    g0541(.A(new_n414), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n223), .A2(new_n497), .A3(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n223), .A2(G179), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n281), .A3(G200), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n744), .A2(new_n372), .B1(new_n344), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n281), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT89), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT89), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(G77), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n223), .A2(new_n497), .A3(new_n369), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n754), .A2(new_n742), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n754), .A2(new_n281), .A3(new_n755), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G50), .A2(new_n757), .B1(new_n758), .B2(G68), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n741), .A2(new_n752), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(G20), .B1(new_n738), .B2(new_n281), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n273), .B1(new_n762), .B2(new_n211), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n761), .A2(G97), .B1(new_n763), .B2(KEYINPUT92), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(KEYINPUT92), .B2(new_n763), .ZN(new_n765));
  INV_X1    g0565(.A(new_n744), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n273), .B1(new_n766), .B2(G322), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n748), .A2(new_n768), .B1(new_n746), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n762), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(G303), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n739), .A2(G329), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n767), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n757), .A2(G326), .B1(new_n761), .B2(G294), .ZN(new_n775));
  INV_X1    g0575(.A(new_n758), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT33), .B(G317), .Z(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n760), .A2(new_n765), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n736), .B1(new_n779), .B2(new_n733), .ZN(new_n780));
  INV_X1    g0580(.A(new_n732), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n641), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n721), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  NAND2_X1  g0584(.A1(new_n630), .A2(new_n638), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n341), .A2(new_n638), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n357), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n355), .B1(new_n348), .B2(KEYINPUT68), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n362), .B1(new_n788), .B2(new_n354), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n789), .B2(new_n786), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n790), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n630), .A3(new_n638), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n722), .B1(new_n794), .B2(new_n705), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n705), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n733), .A2(new_n730), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G77), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n766), .A2(G294), .B1(new_n761), .B2(G97), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G303), .A2(new_n757), .B1(new_n751), .B2(G116), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n404), .B1(new_n762), .B2(new_n344), .C1(new_n211), .C2(new_n746), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G311), .B2(new_n739), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n802), .B(new_n804), .C1(new_n769), .C2(new_n776), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n758), .A2(G150), .B1(new_n766), .B2(G143), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  INV_X1    g0609(.A(new_n751), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n807), .B1(new_n808), .B2(new_n756), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT94), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n273), .B1(new_n746), .B2(new_n373), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G50), .B2(new_n771), .ZN(new_n815));
  INV_X1    g0615(.A(new_n761), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  INV_X1    g0617(.A(new_n739), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n815), .B1(new_n816), .B2(new_n372), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n812), .B2(KEYINPUT94), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n806), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n720), .B(new_n799), .C1(new_n822), .C2(new_n733), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n731), .B2(new_n792), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n796), .A2(new_n824), .ZN(G384));
  OR2_X1    g0625(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(G116), .A4(new_n224), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT36), .Z(new_n829));
  OAI211_X1 g0629(.A(new_n226), .B(G77), .C1(new_n372), .C2(new_n373), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n201), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n255), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n637), .B1(new_n411), .B2(new_n420), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n788), .A2(new_n354), .A3(new_n638), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n793), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n368), .A2(new_n638), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n332), .A2(new_n370), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n607), .B2(new_n597), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n400), .A2(new_n637), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n410), .A2(new_n844), .A3(new_n845), .A4(new_n421), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n386), .A2(G68), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT72), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n395), .A2(new_n381), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n394), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n390), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n253), .B(new_n389), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(new_n399), .B1(new_n407), .B2(new_n408), .ZN(new_n853));
  INV_X1    g0653(.A(new_n637), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n852), .B2(new_n399), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n853), .A2(new_n855), .A3(new_n417), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n846), .B1(new_n856), .B2(new_n845), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n424), .A2(new_n855), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n834), .B1(new_n843), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n410), .A2(new_n844), .A3(new_n421), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(KEYINPUT96), .A3(new_n846), .ZN(new_n866));
  INV_X1    g0666(.A(new_n844), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n424), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT96), .B1(new_n865), .B2(new_n846), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT39), .B1(new_n859), .B2(new_n860), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT97), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT97), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n332), .A2(new_n647), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT95), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n862), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n425), .B1(new_n681), .B2(new_n683), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n610), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n883), .B(new_n885), .Z(new_n886));
  NAND2_X1  g0686(.A1(new_n871), .A2(new_n873), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT98), .B1(new_n695), .B2(new_n638), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT98), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n700), .A2(new_n889), .A3(new_n647), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n890), .A3(new_n685), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n638), .B1(new_n698), .B2(new_n699), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n592), .A2(new_n638), .B1(new_n892), .B2(KEYINPUT31), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n790), .B1(new_n839), .B2(new_n840), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n895), .B(new_n894), .C1(new_n859), .C2(new_n860), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT99), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n425), .A2(new_n894), .ZN(new_n903));
  OAI21_X1  g0703(.A(G330), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n903), .B2(new_n902), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n886), .A2(new_n905), .B1(new_n255), .B2(new_n715), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n886), .A2(new_n905), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n833), .B1(new_n906), .B2(new_n907), .ZN(G367));
  NOR2_X1   g0708(.A1(new_n726), .A2(new_n235), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n734), .B1(new_n219), .B2(new_n333), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n722), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n757), .A2(G143), .B1(new_n761), .B2(G68), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n912), .B1(new_n809), .B2(new_n776), .C1(new_n201), .C2(new_n810), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n818), .A2(new_n808), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n273), .B1(new_n762), .B2(new_n372), .ZN(new_n915));
  INV_X1    g0715(.A(G150), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n744), .A2(new_n916), .B1(new_n276), .B2(new_n746), .ZN(new_n917));
  NOR4_X1   g0717(.A1(new_n913), .A2(new_n914), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(G283), .A2(new_n751), .B1(new_n758), .B2(G294), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n344), .B2(new_n816), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n771), .A2(KEYINPUT46), .A3(G116), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT46), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n762), .B2(new_n489), .ZN(new_n923));
  INV_X1    g0723(.A(G317), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n921), .B(new_n923), .C1(new_n818), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n756), .A2(new_n768), .ZN(new_n926));
  INV_X1    g0726(.A(G303), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n404), .B1(new_n475), .B2(new_n746), .C1(new_n744), .C2(new_n927), .ZN(new_n928));
  NOR4_X1   g0728(.A1(new_n920), .A2(new_n925), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT47), .Z(new_n931));
  AOI21_X1  g0731(.A(new_n911), .B1(new_n931), .B2(new_n733), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n647), .A2(new_n517), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n520), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n624), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n732), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n651), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n647), .A2(new_n676), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n485), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n618), .A2(new_n647), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n943), .B1(new_n649), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n612), .A2(new_n638), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n949), .A2(new_n591), .B1(new_n590), .B2(new_n647), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n485), .A2(new_n944), .B1(new_n618), .B2(new_n647), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT101), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n642), .A2(new_n954), .A3(new_n644), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n649), .A2(new_n947), .A3(KEYINPUT45), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n950), .B2(new_n951), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n953), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n955), .B1(new_n959), .B2(new_n953), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n680), .A2(new_n638), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT29), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n646), .A2(new_n648), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n644), .B2(new_n648), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n642), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n712), .B(new_n965), .C1(new_n644), .C2(new_n648), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n705), .A3(new_n682), .A4(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT102), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n684), .A2(KEYINPUT102), .A3(new_n705), .A4(new_n969), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n962), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n942), .B1(new_n974), .B2(new_n706), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT103), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(KEYINPUT103), .B(new_n942), .C1(new_n974), .C2(new_n706), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n716), .A3(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n947), .A2(KEYINPUT100), .A3(new_n646), .A4(new_n648), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT100), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n965), .B2(new_n951), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n951), .A2(new_n590), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n638), .B1(new_n985), .B2(new_n664), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n937), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n987), .A2(new_n990), .A3(new_n937), .A4(new_n988), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n645), .A2(new_n951), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n979), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT104), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT104), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n979), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n940), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT105), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n717), .B1(new_n975), .B2(new_n976), .ZN(new_n1009));
  AOI211_X1 g0809(.A(KEYINPUT104), .B(new_n1000), .C1(new_n1009), .C2(new_n978), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1004), .B1(new_n979), .B2(new_n1001), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n939), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT105), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(G387));
  NAND2_X1  g0815(.A1(new_n969), .A2(new_n717), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n744), .A2(new_n209), .B1(new_n276), .B2(new_n762), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n748), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(G68), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G159), .A2(new_n757), .B1(new_n758), .B2(new_n245), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n273), .B1(new_n746), .B2(new_n475), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n739), .B2(G150), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n761), .A2(new_n334), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n739), .A2(G326), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n746), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n273), .B1(new_n1026), .B2(G116), .ZN(new_n1027));
  INV_X1    g0827(.A(G294), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n816), .A2(new_n769), .B1(new_n1028), .B2(new_n762), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n757), .A2(G322), .B1(new_n766), .B2(G317), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n927), .B2(new_n810), .C1(new_n768), .C2(new_n776), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1025), .B(new_n1027), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1024), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n733), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n232), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n726), .B1(new_n1040), .B2(G45), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n654), .B1(new_n1041), .B2(new_n723), .ZN(new_n1042));
  XOR2_X1   g0842(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n1043));
  NOR3_X1   g0843(.A1(new_n336), .A2(G50), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n336), .B2(G50), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n266), .C1(new_n373), .C2(new_n276), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1041), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1042), .B(new_n1047), .C1(G107), .C2(new_n219), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n720), .B1(new_n1048), .B2(new_n734), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1039), .B(new_n1049), .C1(new_n644), .C2(new_n781), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n707), .A2(new_n969), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n970), .A2(new_n714), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1016), .B(new_n1050), .C1(new_n1051), .C2(new_n1052), .ZN(G393));
  AND2_X1   g0853(.A1(new_n953), .A2(new_n959), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT107), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n1054), .A2(new_n1055), .A3(new_n645), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1054), .B2(new_n645), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n645), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n716), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n951), .A2(new_n732), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n734), .B1(new_n475), .B2(new_n219), .C1(new_n242), .C2(new_n726), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n722), .A2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n776), .A2(new_n201), .B1(new_n816), .B2(new_n276), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n336), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n751), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n756), .A2(new_n916), .B1(new_n744), .B2(new_n809), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n273), .B1(new_n762), .B2(new_n373), .C1(new_n211), .C2(new_n746), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G143), .B2(new_n739), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n756), .A2(new_n924), .B1(new_n744), .B2(new_n768), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT108), .Z(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n761), .A2(G116), .B1(G294), .B2(new_n1018), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n776), .B2(new_n927), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT109), .Z(new_n1077));
  OAI221_X1 g0877(.A(new_n404), .B1(new_n762), .B2(new_n769), .C1(new_n344), .C2(new_n746), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G322), .B2(new_n739), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1071), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1063), .B1(new_n1081), .B2(new_n733), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1060), .B1(new_n1061), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1059), .A2(new_n970), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n974), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n714), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(G390));
  NAND4_X1  g0887(.A1(new_n841), .A2(G330), .A3(new_n704), .A4(new_n792), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n792), .A2(new_n638), .A3(new_n680), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1088), .A2(new_n1089), .A3(new_n835), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n710), .B1(new_n891), .B2(new_n893), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n841), .B1(new_n1091), .B2(new_n792), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n895), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n792), .A2(new_n704), .A3(G330), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n842), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n793), .A2(new_n835), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1090), .A2(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n425), .A2(new_n1091), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n884), .A2(new_n610), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT110), .Z(new_n1103));
  OAI21_X1  g0903(.A(new_n882), .B1(new_n836), .B2(new_n842), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n874), .A2(new_n878), .A3(new_n875), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n887), .A2(new_n882), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1089), .A2(new_n835), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n841), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1107), .A2(new_n1111), .A3(new_n1088), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n880), .B2(new_n1104), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(new_n1094), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1103), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1112), .B(new_n1102), .C1(new_n1114), .C2(new_n1094), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n714), .A3(new_n1117), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1115), .A2(new_n1113), .A3(new_n716), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n731), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n880), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n722), .B1(new_n245), .B2(new_n798), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n751), .A2(G97), .B1(new_n761), .B2(G77), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n344), .B2(new_n776), .C1(new_n769), .C2(new_n756), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n818), .A2(new_n1028), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n404), .B1(new_n762), .B2(new_n211), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n744), .A2(new_n489), .B1(new_n373), .B2(new_n746), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1129), .A2(KEYINPUT111), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n810), .A2(new_n1131), .B1(new_n1132), .B2(new_n756), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G137), .B2(new_n758), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n771), .A2(G150), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G125), .B2(new_n739), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n273), .B1(new_n201), .B2(new_n746), .C1(new_n744), .C2(new_n817), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G159), .B2(new_n761), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1129), .A2(KEYINPUT111), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1130), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1122), .B1(new_n1142), .B2(new_n733), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1119), .B1(new_n1121), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1118), .A2(new_n1144), .ZN(G378));
  OAI211_X1 g0945(.A(G330), .B(new_n896), .C1(new_n900), .C2(new_n901), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n883), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n862), .C1(new_n882), .C2(new_n880), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n596), .A2(new_n359), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n261), .A2(new_n637), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT55), .Z(new_n1152));
  XNOR2_X1  g0952(.A(new_n1150), .B(new_n1152), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT113), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1148), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1155), .A2(new_n731), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n720), .B1(new_n201), .B2(new_n797), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT112), .Z(new_n1161));
  OAI22_X1  g0961(.A1(new_n776), .A2(new_n817), .B1(new_n816), .B2(new_n916), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n766), .A2(G128), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1131), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n771), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1018), .A2(G137), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1162), .B(new_n1167), .C1(G125), .C2(new_n757), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n263), .B(new_n264), .C1(new_n746), .C2(new_n809), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n739), .B2(G124), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n758), .A2(G97), .B1(new_n761), .B2(G68), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n489), .B2(new_n756), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n273), .A2(G41), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n276), .B2(new_n762), .C1(new_n818), .C2(new_n769), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n766), .A2(G107), .B1(G58), .B2(new_n1026), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n333), .B2(new_n748), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1177), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n209), .C1(G33), .C2(G41), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1174), .A2(new_n1182), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1161), .B1(new_n1186), .B2(new_n733), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1158), .A2(new_n717), .B1(new_n1159), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT114), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n884), .A2(new_n610), .A3(new_n1100), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1117), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1117), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1158), .B(KEYINPUT57), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n714), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1117), .A2(new_n1190), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT114), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1117), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1158), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1188), .B1(new_n1194), .B2(new_n1199), .ZN(G375));
  AOI22_X1  g1000(.A1(new_n1091), .A2(new_n895), .B1(new_n1095), .B2(new_n842), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1088), .A2(new_n1089), .A3(new_n835), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1201), .A2(new_n836), .B1(new_n1202), .B2(new_n1092), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1103), .B(new_n942), .C1(new_n1190), .C2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n842), .A2(new_n730), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n722), .B1(G68), .B2(new_n798), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n748), .A2(new_n916), .B1(new_n762), .B2(new_n809), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n273), .B1(new_n372), .B2(new_n746), .C1(new_n818), .C2(new_n1132), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G137), .C2(new_n766), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n756), .A2(new_n817), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT117), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n758), .A2(new_n1164), .B1(new_n761), .B2(G50), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G294), .A2(new_n757), .B1(new_n758), .B2(G116), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n344), .B2(new_n810), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT115), .Z(new_n1216));
  AOI22_X1  g1016(.A1(new_n739), .A2(G303), .B1(G97), .B2(new_n771), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT116), .Z(new_n1218));
  OAI21_X1  g1018(.A(new_n404), .B1(new_n746), .B2(new_n276), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n766), .B2(G283), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1023), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1213), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1206), .B1(new_n1222), .B2(new_n733), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1203), .A2(new_n717), .B1(new_n1205), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1204), .A2(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT118), .Z(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1014), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(G375), .ZN(G407));
  INV_X1    g1031(.A(G343), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G213), .ZN(new_n1233));
  OR3_X1    g1033(.A1(G375), .A2(G378), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1008), .A2(new_n1013), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(new_n783), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT122), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1006), .B2(G390), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1012), .A2(new_n1245), .A3(new_n1237), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G390), .B(new_n939), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1012), .B2(new_n1237), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1242), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n1242), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1244), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1236), .B1(new_n1254), .B2(KEYINPUT61), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1253), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT123), .B1(new_n1006), .B2(G390), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1252), .B1(new_n1259), .B2(new_n1242), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1256), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(KEYINPUT126), .A3(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G378), .B(new_n1188), .C1(new_n1194), .C2(new_n1199), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1198), .A2(new_n942), .A3(new_n1158), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1188), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1228), .A2(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1264), .A2(new_n1267), .B1(G213), .B2(new_n1232), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1190), .B2(new_n1203), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n651), .B1(new_n1190), .B2(new_n1203), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1101), .A3(new_n1275), .A4(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT119), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT119), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1099), .A2(new_n1278), .A3(KEYINPUT60), .A4(new_n1101), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1224), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1224), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(new_n1273), .C2(new_n1280), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1268), .A2(new_n1286), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1232), .A2(G213), .A3(G2897), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT120), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT121), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1272), .B1(new_n1279), .B2(new_n1277), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1283), .B1(new_n1293), .B2(new_n1284), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1281), .A2(G384), .A3(new_n1224), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(KEYINPUT120), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1290), .B(KEYINPUT121), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1291), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT121), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1289), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1296), .B2(KEYINPUT120), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1296), .A2(KEYINPUT120), .A3(new_n1292), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1233), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1288), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1255), .A2(new_n1263), .A3(new_n1287), .A4(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1306), .A2(new_n1311), .A3(new_n1233), .A4(new_n1286), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(new_n1262), .C1(new_n1268), .C2(new_n1305), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1268), .B2(new_n1286), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1254), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(G375), .A2(new_n1228), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1264), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1286), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1317), .B(new_n1264), .C1(KEYINPUT127), .C2(new_n1296), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1254), .ZN(G402));
endmodule


