//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT65), .B(G244), .ZN(new_n212));
  AND2_X1   g0012(.A1(new_n212), .A2(G77), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n208), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n202), .A2(new_n203), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR4_X1   g0028(.A1(new_n211), .A2(new_n222), .A3(new_n223), .A4(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  INV_X1    g0031(.A(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  INV_X1    g0039(.A(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n203), .A2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n226), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n249), .B1(new_n250), .B2(new_n251), .C1(new_n253), .C2(new_n201), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n227), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n257), .A2(KEYINPUT11), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(KEYINPUT11), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT12), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n260), .A2(new_n261), .A3(G1), .ZN(new_n264));
  INV_X1    g0064(.A(new_n249), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n260), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n258), .A2(new_n259), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n255), .A2(new_n227), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n261), .A2(new_n226), .A3(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT71), .B1(new_n271), .B2(new_n256), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n203), .B1(new_n276), .B2(KEYINPUT12), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI211_X1 g0082(.A(G232), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G97), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n232), .B1(new_n288), .B2(new_n289), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n280), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n280), .A3(G274), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(KEYINPUT73), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT73), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  INV_X1    g0105(.A(new_n227), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n279), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n307), .B2(new_n301), .ZN(new_n308));
  INV_X1    g0108(.A(G238), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n280), .A2(new_n310), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n303), .A2(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT13), .B1(new_n298), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n302), .A2(KEYINPUT73), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n307), .A2(new_n304), .A3(new_n301), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n301), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n315), .A2(new_n316), .B1(G238), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(G226), .B(new_n296), .C1(new_n281), .C2(new_n282), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n287), .B2(new_n293), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n285), .B2(new_n291), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n314), .B(new_n319), .C1(new_n322), .C2(new_n280), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n313), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n278), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n313), .A2(new_n323), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n327), .A2(new_n331), .A3(G169), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n313), .A2(new_n323), .A3(G179), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n327), .B2(G169), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT74), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT14), .B1(new_n324), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(new_n333), .A4(new_n332), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n278), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n330), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT8), .B(G58), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n275), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n268), .A2(new_n263), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n346), .A2(new_n347), .B1(new_n263), .B2(new_n345), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT77), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n288), .A2(new_n226), .A3(new_n289), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n289), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT76), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  OAI21_X1  g0156(.A(G68), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n226), .B1(new_n224), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n252), .A2(G159), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT16), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n281), .A2(new_n282), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT7), .B1(new_n364), .B2(new_n226), .ZN(new_n365));
  INV_X1    g0165(.A(new_n354), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT75), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n359), .B2(new_n361), .ZN(new_n369));
  INV_X1    g0169(.A(new_n359), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n360), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n256), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n349), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n349), .B(KEYINPUT78), .C1(new_n363), .C2(new_n373), .ZN(new_n377));
  OAI211_X1 g0177(.A(G223), .B(new_n296), .C1(new_n281), .C2(new_n282), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT79), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n295), .A2(G1698), .B1(G33), .B2(G87), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n280), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n280), .A2(G232), .A3(new_n310), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n302), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n386), .B(KEYINPUT80), .ZN(new_n387));
  OAI21_X1  g0187(.A(G169), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT80), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n386), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n290), .A2(G226), .ZN(new_n392));
  INV_X1    g0192(.A(G87), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n392), .A2(new_n296), .B1(new_n287), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n381), .B2(new_n380), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(new_n280), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n388), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n376), .A2(new_n377), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  OAI21_X1  g0200(.A(G200), .B1(new_n384), .B2(new_n387), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n391), .B(G190), .C1(new_n395), .C2(new_n280), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT77), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n348), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n357), .A2(new_n362), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n372), .A2(new_n256), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n403), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n401), .A2(new_n402), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT17), .B1(new_n413), .B2(new_n374), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n398), .A2(new_n400), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n376), .A2(new_n397), .A3(new_n377), .A4(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n302), .B1(new_n232), .B2(new_n311), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n364), .A2(G1698), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(G222), .B1(G77), .B2(new_n364), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT68), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n364), .B2(new_n296), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n290), .A2(KEYINPUT68), .A3(G1698), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(G223), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT69), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n280), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT69), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G190), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G150), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n344), .A2(new_n250), .B1(new_n432), .B2(new_n253), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(G20), .B2(new_n204), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n268), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n275), .A2(G50), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n347), .A2(new_n436), .B1(G50), .B2(new_n263), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT9), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n437), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT9), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n434), .C2(new_n268), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n429), .B2(new_n325), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT10), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n429), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G200), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT10), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n430), .A4(new_n442), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n445), .A2(new_n337), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n435), .A2(new_n437), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n429), .B2(new_n389), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n318), .A2(new_n212), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n302), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT70), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT70), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n457), .A3(new_n302), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n420), .A2(G232), .B1(G107), .B2(new_n364), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n423), .A2(G238), .A3(new_n424), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n280), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n337), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n462), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n389), .A3(new_n456), .A4(new_n458), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n273), .A2(G77), .A3(new_n275), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n271), .A2(new_n251), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G20), .A2(G77), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT15), .B(G87), .ZN(new_n469));
  OAI221_X1 g0269(.A(new_n468), .B1(new_n344), .B2(new_n253), .C1(new_n250), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n256), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n463), .A2(new_n465), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n464), .A2(new_n456), .A3(new_n458), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  INV_X1    g0275(.A(new_n472), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n476), .C1(new_n474), .C2(new_n328), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n453), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n343), .A2(new_n418), .A3(new_n449), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT83), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G41), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n299), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n300), .A2(G1), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n307), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G270), .A3(new_n280), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(G264), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT86), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n290), .A2(KEYINPUT86), .A3(G264), .A4(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G257), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n288), .B2(new_n289), .ZN(new_n500));
  XOR2_X1   g0300(.A(KEYINPUT87), .B(G303), .Z(new_n501));
  AOI22_X1  g0301(.A1(new_n296), .A2(new_n500), .B1(new_n501), .B2(new_n364), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n493), .B1(new_n503), .B2(new_n280), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n504), .A2(new_n328), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n243), .B1(new_n274), .B2(G33), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n270), .A2(new_n272), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n271), .A2(new_n243), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n243), .A2(G20), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n256), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n226), .C1(G33), .C2(new_n293), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT20), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AND4_X1   g0313(.A1(KEYINPUT20), .A2(new_n512), .A3(new_n256), .A4(new_n509), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n507), .B(new_n508), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n504), .B2(G200), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n504), .A2(KEYINPUT21), .A3(G169), .A4(new_n515), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n280), .B1(new_n498), .B2(new_n502), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n515), .B(G169), .C1(new_n519), .C2(new_n492), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n519), .A2(new_n492), .A3(new_n389), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n515), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n274), .B(G45), .C1(new_n299), .C2(KEYINPUT5), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n482), .A2(G41), .ZN(new_n528));
  OAI211_X1 g0328(.A(G257), .B(new_n280), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n490), .A2(KEYINPUT84), .A3(G257), .A4(new_n280), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n317), .A2(new_n527), .A3(new_n305), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n531), .A2(new_n532), .B1(new_n485), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(new_n296), .C1(new_n281), .C2(new_n282), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n511), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT82), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(new_n541), .A3(new_n537), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n534), .B1(new_n543), .B2(new_n280), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n337), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n534), .B(new_n389), .C1(new_n543), .C2(new_n280), .ZN(new_n546));
  OAI21_X1  g0346(.A(G107), .B1(new_n355), .B2(new_n356), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n293), .A2(new_n240), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n240), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n268), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n263), .A2(G97), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n347), .B1(new_n274), .B2(G33), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(G97), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n546), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n544), .A2(KEYINPUT85), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n536), .A2(new_n537), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n535), .A2(new_n511), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n536), .A2(new_n541), .A3(new_n537), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n541), .B1(new_n536), .B2(new_n537), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n317), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT85), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n534), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(new_n570), .A3(G200), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT76), .B1(new_n365), .B2(new_n366), .ZN(new_n572));
  INV_X1    g0372(.A(new_n356), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n240), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n554), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n256), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n534), .B(G190), .C1(new_n543), .C2(new_n280), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n576), .A2(new_n577), .A3(new_n558), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n545), .A2(new_n561), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n580));
  OAI211_X1 g0380(.A(G250), .B(new_n296), .C1(new_n281), .C2(new_n282), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G294), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n317), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT88), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT88), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n586), .A3(new_n317), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n490), .A2(G264), .A3(new_n280), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n488), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n584), .A2(new_n488), .A3(new_n588), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n592), .A2(new_n389), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n226), .B(G87), .C1(new_n281), .C2(new_n282), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT22), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT22), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n290), .A2(new_n597), .A3(new_n226), .A4(G87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G116), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(G20), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT23), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n226), .B2(G107), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n240), .A2(KEYINPUT23), .A3(G20), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n600), .B1(new_n599), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n256), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n271), .A2(new_n240), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT25), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(G107), .B2(new_n557), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n594), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n469), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n557), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n290), .A2(new_n226), .A3(G68), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n393), .A2(new_n293), .A3(new_n240), .ZN(new_n618));
  OAI211_X1 g0418(.A(KEYINPUT19), .B(new_n618), .C1(new_n294), .C2(G20), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n250), .A2(new_n293), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n617), .B(new_n619), .C1(KEYINPUT19), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n256), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n469), .A2(new_n271), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n616), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n309), .A2(new_n296), .ZN(new_n625));
  INV_X1    g0425(.A(G244), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G1698), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n625), .B(new_n627), .C1(new_n281), .C2(new_n282), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n280), .B1(new_n628), .B2(new_n601), .ZN(new_n629));
  INV_X1    g0429(.A(G250), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n300), .B2(G1), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n274), .A2(new_n305), .A3(G45), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n280), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n337), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n601), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n317), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n389), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n624), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n621), .A2(new_n256), .B1(new_n271), .B2(new_n469), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n557), .A2(G87), .ZN(new_n640));
  OAI21_X1  g0440(.A(G200), .B1(new_n629), .B2(new_n633), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(G190), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n592), .A2(new_n325), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n590), .B2(G190), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n609), .A3(new_n612), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n614), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n480), .A2(new_n526), .A3(new_n579), .A4(new_n648), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n412), .A2(new_n414), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n278), .B1(new_n336), .B2(new_n340), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n473), .A2(KEYINPUT91), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT91), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n463), .A2(new_n465), .A3(new_n653), .A4(new_n472), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n330), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n650), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n397), .A2(new_n374), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(new_n399), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n444), .A2(new_n448), .A3(KEYINPUT92), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT92), .B1(new_n444), .B2(new_n448), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n660), .A2(new_n663), .B1(new_n450), .B2(new_n452), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n638), .B(KEYINPUT89), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n576), .A2(new_n558), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n545), .A3(new_n546), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n638), .A2(new_n643), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT90), .ZN(new_n673));
  AOI21_X1  g0473(.A(G169), .B1(new_n568), .B2(new_n534), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n560), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n667), .A2(KEYINPUT90), .A3(new_n545), .A4(new_n546), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n571), .A2(new_n578), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n668), .A3(new_n647), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n591), .A2(new_n593), .B1(new_n609), .B2(new_n612), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n525), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n672), .B1(new_n682), .B2(new_n644), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n664), .B1(new_n479), .B2(new_n683), .ZN(G369));
  NAND2_X1  g0484(.A1(new_n262), .A2(new_n226), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n680), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT93), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n613), .A2(new_n690), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n614), .A2(new_n647), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n515), .A2(new_n690), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n525), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n517), .A2(new_n525), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n690), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n525), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n692), .B2(new_n694), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n614), .A2(new_n690), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n209), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  NOR4_X1   g0511(.A1(new_n711), .A2(new_n274), .A3(G116), .A4(new_n618), .ZN(new_n712));
  INV_X1    g0512(.A(new_n225), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n711), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  NOR3_X1   g0515(.A1(new_n683), .A2(KEYINPUT29), .A3(new_n690), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n671), .B1(new_n668), .B2(new_n669), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n665), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n614), .A2(new_n522), .A3(new_n524), .A4(new_n518), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n579), .A2(new_n720), .A3(new_n644), .A4(new_n647), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n690), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n636), .A2(new_n584), .A3(new_n588), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n568), .A2(new_n728), .A3(new_n534), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n493), .B(G179), .C1(new_n503), .C2(new_n280), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n531), .A2(new_n532), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n488), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n317), .B2(new_n567), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(KEYINPUT30), .A3(new_n523), .A4(new_n728), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n636), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n504), .A2(new_n544), .A3(new_n592), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n731), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT31), .B1(new_n738), .B2(new_n690), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n526), .A2(new_n648), .A3(new_n579), .A4(new_n704), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n726), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n725), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n715), .B1(new_n746), .B2(G1), .ZN(G364));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n227), .B1(G20), .B2(new_n337), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n710), .A2(new_n290), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n225), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(G45), .B2(new_n247), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n209), .A2(new_n290), .ZN(new_n756));
  XOR2_X1   g0556(.A(G355), .B(KEYINPUT94), .Z(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n209), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n752), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n261), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n274), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n711), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n226), .A2(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n393), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n226), .A2(new_n389), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n328), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n226), .B1(new_n772), .B2(G190), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n201), .B1(new_n773), .B2(new_n293), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n769), .A2(G190), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n767), .B(new_n774), .C1(G68), .C2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n765), .A2(new_n328), .A3(G200), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n290), .B1(new_n777), .B2(new_n240), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n768), .B(KEYINPUT95), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n778), .B1(new_n782), .B2(G77), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n772), .A2(G20), .A3(new_n328), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT32), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OR3_X1    g0589(.A1(new_n787), .A2(KEYINPUT32), .A3(new_n788), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n776), .A2(new_n783), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n328), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n202), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G311), .A2(new_n782), .B1(new_n794), .B2(G322), .ZN(new_n800));
  INV_X1    g0600(.A(new_n787), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G329), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(KEYINPUT100), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT100), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n775), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n800), .B(new_n802), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n364), .B1(new_n766), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT99), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT99), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT98), .B(G326), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n770), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n777), .ZN(new_n815));
  INV_X1    g0615(.A(new_n773), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(G283), .B1(new_n816), .B2(G294), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n791), .A2(new_n799), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n764), .B1(new_n819), .B2(new_n751), .ZN(new_n820));
  INV_X1    g0620(.A(new_n750), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n700), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n763), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n701), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n700), .A2(G330), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n682), .A2(new_n644), .ZN(new_n827));
  INV_X1    g0627(.A(new_n672), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n690), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n476), .A2(new_n704), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n477), .A2(new_n473), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n652), .A2(new_n654), .A3(new_n830), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n829), .B(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n763), .B1(new_n836), .B2(new_n744), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n744), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n751), .A2(new_n748), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n763), .B1(G77), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G116), .A2(new_n782), .B1(new_n794), .B2(G294), .ZN(new_n842));
  INV_X1    g0642(.A(new_n775), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n843), .A2(new_n844), .B1(new_n771), .B2(new_n809), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n777), .A2(new_n393), .B1(new_n766), .B2(new_n240), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n801), .A2(G311), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n290), .B1(new_n816), .B2(G97), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n842), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n775), .A2(G150), .B1(new_n770), .B2(G137), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n781), .B2(new_n788), .ZN(new_n852));
  INV_X1    g0652(.A(new_n798), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(G143), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n290), .B1(new_n773), .B2(new_n202), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n777), .A2(new_n203), .B1(new_n766), .B2(new_n201), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n801), .C2(G132), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n850), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n841), .B1(new_n861), .B2(new_n751), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n749), .B2(new_n835), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n838), .A2(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n760), .A2(new_n274), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n834), .B1(new_n741), .B2(new_n742), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n342), .A2(new_n690), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n651), .A2(new_n330), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n336), .B2(new_n340), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n688), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n376), .A2(new_n377), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT37), .B1(new_n403), .B2(new_n410), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n398), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT102), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT102), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n398), .A2(new_n873), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n367), .A2(KEYINPUT101), .A3(new_n369), .A4(new_n371), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n883), .A2(new_n407), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n349), .B1(new_n885), .B2(new_n373), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n886), .A2(new_n397), .B1(new_n403), .B2(new_n410), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n872), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n415), .B2(new_n417), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n889), .B1(new_n876), .B2(new_n878), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n892), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n871), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT103), .B1(new_n898), .B2(KEYINPUT40), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n870), .B1(new_n343), .B2(new_n867), .ZN(new_n900));
  INV_X1    g0700(.A(new_n740), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n742), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n835), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n891), .B2(new_n893), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n896), .A2(new_n895), .A3(new_n892), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT103), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n899), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n873), .B(new_n658), .C1(new_n374), .C2(new_n413), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n879), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n873), .B1(new_n659), .B2(new_n650), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n907), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n866), .B(KEYINPUT40), .C1(new_n869), .C2(new_n870), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n912), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT104), .Z(new_n922));
  NAND2_X1  g0722(.A1(new_n480), .A2(new_n903), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n726), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n922), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n906), .A2(new_n907), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n473), .A2(new_n690), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n829), .B2(new_n835), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(new_n900), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n927), .A2(new_n930), .B1(new_n659), .B2(new_n872), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n651), .A2(new_n704), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT39), .B1(new_n906), .B2(new_n907), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n876), .A2(new_n878), .B1(new_n913), .B2(KEYINPUT37), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n895), .B1(new_n934), .B2(new_n916), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n894), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n932), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n660), .A2(new_n663), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n453), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n719), .A2(new_n721), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT29), .B1(new_n942), .B2(new_n690), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n579), .A2(new_n647), .A3(new_n720), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n669), .B1(new_n944), .B2(new_n677), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n723), .B(new_n704), .C1(new_n945), .C2(new_n672), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n479), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n939), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n865), .B1(new_n926), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n926), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n227), .A2(new_n226), .A3(new_n243), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT36), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n713), .A2(G77), .A3(new_n358), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(G50), .B2(new_n203), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(G1), .A3(new_n261), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n951), .A2(new_n956), .A3(new_n959), .ZN(G367));
  NAND2_X1  g0760(.A1(new_n639), .A2(new_n640), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n690), .ZN(new_n962));
  MUX2_X1   g0762(.A(new_n666), .B(new_n669), .S(new_n962), .Z(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n667), .A2(new_n690), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n579), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n561), .A2(new_n545), .A3(new_n690), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n706), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n970), .A2(KEYINPUT42), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n579), .A2(new_n680), .A3(new_n966), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n690), .B1(new_n972), .B2(new_n668), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n970), .B2(KEYINPUT42), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n965), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n963), .A2(new_n964), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n969), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n703), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n711), .B(KEYINPUT41), .Z(new_n981));
  OR3_X1    g0781(.A1(new_n708), .A2(KEYINPUT44), .A3(new_n969), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT44), .B1(new_n708), .B2(new_n969), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT45), .B1(new_n708), .B2(new_n969), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n703), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(KEYINPUT105), .A3(new_n702), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n701), .A2(new_n706), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n705), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT106), .B1(new_n695), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n701), .A2(new_n706), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n994), .B1(new_n991), .B2(new_n995), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n988), .A2(new_n746), .A3(new_n989), .A4(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n981), .B1(new_n999), .B2(new_n746), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n980), .B1(new_n1000), .B2(new_n762), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n753), .A2(new_n237), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n752), .B1(new_n209), .B2(new_n469), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n763), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n963), .B2(new_n750), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n766), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(G116), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT46), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n770), .A2(G311), .B1(G107), .B2(new_n816), .ZN(new_n1009));
  INV_X1    g0809(.A(G294), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1009), .C1(new_n1010), .C2(new_n843), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n777), .A2(new_n293), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n290), .B(new_n1012), .C1(new_n801), .C2(G317), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n844), .B2(new_n781), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1011), .B(new_n1014), .C1(new_n853), .C2(new_n501), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n816), .A2(G68), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n793), .B2(new_n432), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n770), .A2(G143), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n202), .B2(new_n766), .C1(new_n843), .C2(new_n788), .ZN(new_n1020));
  INV_X1    g0820(.A(G137), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n781), .A2(new_n201), .B1(new_n787), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n290), .B1(new_n777), .B2(new_n251), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT108), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1015), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT109), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n751), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1005), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1001), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n998), .A2(new_n762), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n775), .A2(G311), .B1(new_n770), .B2(G322), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n501), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n781), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n853), .B2(G317), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT48), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(KEYINPUT48), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1006), .A2(G294), .B1(new_n816), .B2(G283), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT49), .Z(new_n1041));
  AND2_X1   g0841(.A1(new_n801), .A2(new_n813), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n364), .B1(new_n777), .B2(new_n243), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n364), .B(new_n1012), .C1(new_n794), .C2(G50), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n203), .B2(new_n781), .C1(new_n432), .C2(new_n787), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n816), .A2(new_n615), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n771), .B2(new_n788), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n843), .A2(new_n344), .B1(new_n251), .B2(new_n766), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n751), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n234), .A2(G45), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT110), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n345), .A2(new_n201), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT50), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n618), .A2(G116), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n300), .C1(new_n203), .C2(new_n251), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1053), .B(new_n753), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(G107), .B2(new_n209), .C1(new_n1056), .C2(new_n756), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n823), .B1(new_n1059), .B2(new_n752), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1051), .B(new_n1060), .C1(new_n695), .C2(new_n821), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n998), .A2(new_n746), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n711), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n998), .A2(new_n746), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1032), .B(new_n1061), .C1(new_n1063), .C2(new_n1064), .ZN(G393));
  NOR2_X1   g0865(.A1(new_n969), .A2(new_n821), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT111), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n794), .A2(G311), .B1(G317), .B2(new_n770), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n364), .B1(new_n240), .B2(new_n777), .C1(new_n781), .C2(new_n1010), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G322), .B2(new_n801), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n843), .A2(new_n1034), .B1(new_n844), .B2(new_n766), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G116), .B2(new_n816), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n793), .A2(new_n788), .B1(new_n432), .B2(new_n771), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n290), .B1(new_n393), .B2(new_n777), .C1(new_n781), .C2(new_n344), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G143), .B2(new_n801), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n773), .A2(new_n251), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n766), .A2(new_n203), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(G50), .C2(new_n775), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1076), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1029), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n244), .A2(new_n710), .A3(new_n290), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n752), .B1(new_n209), .B2(new_n293), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n763), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OR3_X1    g0886(.A1(new_n1067), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n986), .B(new_n702), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n761), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n711), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1088), .B2(new_n1062), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(new_n999), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G390));
  OAI21_X1  g0893(.A(new_n932), .B1(new_n929), .B2(new_n900), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n933), .A3(new_n937), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n743), .B(new_n835), .C1(new_n869), .C2(new_n870), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n894), .A2(new_n935), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n928), .B1(new_n722), .B2(new_n835), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n932), .C1(new_n900), .C2(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1095), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n480), .A2(new_n743), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n903), .A2(G330), .A3(new_n835), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n900), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n929), .B1(new_n1096), .B2(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1104), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n948), .B(new_n1102), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1100), .A2(new_n1101), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT112), .B1(new_n1108), .B2(new_n1090), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1101), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1107), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1095), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT112), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n711), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1110), .A2(new_n762), .A3(new_n1112), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n933), .A2(new_n748), .A3(new_n937), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n840), .A2(new_n345), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n775), .A2(G137), .B1(G159), .B2(new_n816), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n771), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n782), .A2(new_n1125), .B1(new_n801), .B2(G125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n290), .B1(new_n777), .B2(new_n201), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n794), .B2(G132), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT53), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n766), .B2(new_n432), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1006), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1123), .B(new_n1129), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT113), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n843), .A2(new_n240), .B1(new_n771), .B2(new_n844), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1079), .B(new_n1137), .C1(G68), .C2(new_n815), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n290), .B(new_n767), .C1(new_n782), .C2(G97), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n801), .A2(G294), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n794), .A2(G116), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1135), .A2(new_n1136), .A3(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n823), .B(new_n1120), .C1(new_n1143), .C2(new_n751), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1118), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1117), .A2(new_n1147), .ZN(G378));
  INV_X1    g0948(.A(new_n939), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n453), .B1(new_n661), .B2(new_n662), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n872), .B1(new_n435), .B2(new_n437), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT116), .Z(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1152), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n453), .B(new_n1155), .C1(new_n661), .C2(new_n662), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1154), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(G330), .B1(new_n919), .B2(new_n920), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n911), .C2(new_n899), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1159), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n920), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n726), .B1(new_n1097), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n912), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1149), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n898), .A2(KEYINPUT103), .A3(KEYINPUT40), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1159), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n912), .A2(new_n1164), .A3(new_n1162), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n939), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n480), .B1(new_n716), .B2(new_n724), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n664), .A3(new_n1102), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1166), .A2(new_n1172), .B1(new_n1175), .B2(new_n1113), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n711), .B1(new_n1176), .B2(KEYINPUT57), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1113), .A2(new_n1175), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1178), .A2(KEYINPUT57), .A3(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1159), .A2(new_n748), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n763), .B1(G50), .B2(new_n840), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G50), .B1(new_n289), .B2(new_n299), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n775), .A2(G97), .B1(new_n815), .B2(G58), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n1016), .C1(new_n243), .C2(new_n771), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G41), .B(new_n290), .C1(new_n1006), .C2(G77), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(KEYINPUT114), .B2(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n781), .A2(new_n469), .B1(new_n787), .B2(new_n844), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G107), .B2(new_n794), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(KEYINPUT114), .C2(new_n1187), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n801), .A2(G124), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n815), .C2(G159), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n770), .A2(G125), .B1(G150), .B2(new_n816), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT115), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n775), .A2(G132), .B1(new_n1006), .B2(new_n1125), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n793), .B2(new_n1122), .C1(new_n1021), .C2(new_n781), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT59), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1194), .B(new_n1195), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1200), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1193), .B1(new_n1192), .B2(new_n1191), .C1(new_n1202), .C2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1183), .B1(new_n1205), .B2(new_n751), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1178), .A2(new_n762), .B1(new_n1182), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(G375));
  INV_X1    g1008(.A(new_n981), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1104), .A2(new_n1096), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n929), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1104), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1174), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1107), .A2(new_n1209), .A3(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT117), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1047), .B1(new_n771), .B2(new_n1010), .C1(new_n793), .C2(new_n844), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n781), .A2(new_n240), .B1(new_n243), .B2(new_n843), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(KEYINPUT118), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n364), .B1(new_n777), .B2(new_n251), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT119), .Z(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(KEYINPUT118), .C2(new_n1218), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n787), .A2(new_n809), .B1(new_n293), .B2(new_n766), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT120), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n781), .A2(new_n432), .B1(new_n201), .B2(new_n773), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT122), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n843), .A2(new_n1124), .B1(new_n788), .B2(new_n766), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n290), .B1(new_n202), .B2(new_n777), .C1(new_n787), .C2(new_n1122), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(G132), .C2(new_n770), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n798), .B2(new_n1021), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1227), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n751), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n763), .C1(G68), .C2(new_n840), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n900), .B2(new_n748), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1239), .B2(new_n762), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1216), .A2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT123), .Z(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(G381));
  INV_X1    g1043(.A(new_n1116), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1113), .A2(new_n711), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(KEYINPUT112), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1146), .B1(new_n1246), .B2(new_n1115), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1181), .A2(new_n1247), .A3(new_n1207), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1001), .A2(new_n1030), .A3(new_n1092), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1250), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1242), .A3(new_n1251), .ZN(G407));
  NAND2_X1  g1052(.A1(new_n689), .A2(G213), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT124), .Z(new_n1254));
  NAND2_X1  g1054(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  OAI211_X1 g1056(.A(G378), .B(new_n1207), .C1(new_n1177), .C2(new_n1180), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1178), .A2(new_n1209), .A3(new_n1179), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1207), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1247), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1214), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n711), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1107), .B2(new_n1214), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1240), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G384), .B(new_n1240), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1261), .A2(new_n1253), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n689), .A2(G213), .A3(G2897), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1268), .A2(new_n1269), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT125), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1268), .A2(new_n1279), .A3(new_n1269), .A4(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1254), .A2(G2897), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1275), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  AOI211_X1 g1085(.A(KEYINPUT126), .B(new_n1283), .C1(new_n1278), .C2(new_n1280), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1261), .A2(new_n1253), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1254), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1250), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(G393), .B(G396), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1092), .B1(new_n1001), .B2(new_n1030), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1292), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(G390), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1293), .B1(new_n1297), .B2(new_n1250), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1296), .A2(new_n1298), .A3(KEYINPUT61), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1274), .A2(new_n1289), .A3(new_n1291), .A4(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1290), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1272), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1290), .A2(KEYINPUT62), .A3(new_n1271), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1300), .B1(new_n1307), .B2(new_n1308), .ZN(G405));
  OAI211_X1 g1109(.A(KEYINPUT127), .B(new_n1270), .C1(new_n1296), .C2(new_n1298), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1294), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1297), .A2(new_n1250), .A3(new_n1293), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1270), .A2(KEYINPUT127), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1257), .B1(KEYINPUT127), .B2(new_n1270), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n1247), .B2(G375), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1315), .B(new_n1317), .ZN(G402));
endmodule


