//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n465), .A2(new_n462), .A3(G101), .A4(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n462), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n475), .B2(new_n462), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n472), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n471), .B1(new_n476), .B2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n468), .A2(new_n469), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n486), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(G136), .B2(new_n494), .ZN(G162));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(G2104), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n468), .B2(new_n469), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n504), .B(new_n506), .C1(new_n469), .C2(new_n468), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n504), .B1(new_n468), .B2(new_n469), .ZN(new_n508));
  INV_X1    g083(.A(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n507), .B2(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT6), .B(G651), .Z(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n515), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  XNOR2_X1  g095(.A(new_n512), .B(KEYINPUT71), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(new_n512), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n517), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT6), .B(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(G543), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n514), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n534), .A2(G52), .B1(G90), .B2(new_n526), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n534), .A2(G43), .B1(G81), .B2(new_n526), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND4_X1  g128(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n532), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n525), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G299));
  NAND2_X1  g135(.A1(new_n534), .A2(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n562));
  INV_X1    g137(.A(G87), .ZN(new_n563));
  INV_X1    g138(.A(new_n526), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT74), .ZN(G288));
  NAND2_X1  g141(.A1(new_n512), .A2(G86), .ZN(new_n567));
  NAND2_X1  g142(.A1(G48), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n517), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(G73), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n512), .B2(G61), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n514), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n569), .B1(new_n572), .B2(KEYINPUT75), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n514), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G305));
  NAND2_X1  g150(.A1(new_n521), .A2(G60), .ZN(new_n576));
  NAND2_X1  g151(.A1(G72), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n514), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(G85), .ZN(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n533), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(G54), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n533), .A2(new_n585), .B1(new_n514), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT76), .Z(new_n588));
  NAND2_X1  g163(.A1(new_n526), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G321));
  MUX2_X1   g169(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g170(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n592), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n592), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n487), .A2(G123), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n462), .A2(G111), .ZN(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G135), .B2(new_n494), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT81), .Z(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2096), .Z(new_n609));
  INV_X1    g184(.A(G2104), .ZN(new_n610));
  NOR3_X1   g185(.A1(new_n482), .A2(new_n610), .A3(G2105), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT79), .B(G2100), .ZN(new_n618));
  OAI22_X1  g193(.A1(new_n614), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n616), .B2(new_n614), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n617), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n609), .A2(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n628), .B(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT83), .Z(G401));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G1981), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1986), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G23), .ZN(new_n676));
  INV_X1    g251(.A(new_n565), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n675), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT33), .B(G1976), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n675), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1971), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  AND2_X1   g260(.A1(new_n675), .A2(G6), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G305), .B2(G16), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n678), .A2(new_n679), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n684), .B(new_n688), .C1(new_n685), .C2(new_n687), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(KEYINPUT34), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(KEYINPUT34), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT85), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT85), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n487), .A2(G119), .ZN(new_n697));
  OR2_X1    g272(.A1(G95), .A2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n698), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G131), .B2(new_n494), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n696), .B1(new_n701), .B2(new_n695), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n675), .A2(G24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n582), .B2(new_n675), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  OR4_X1    g282(.A1(new_n690), .A2(new_n691), .A3(new_n704), .A4(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n494), .A2(G141), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n487), .A2(G129), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT26), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n610), .A2(G2105), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n717), .A2(new_n718), .B1(G105), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n713), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(new_n692), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n692), .B2(G32), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1341), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n547), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G19), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G34), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(G34), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n695), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G160), .B2(G29), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(G2084), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(G2084), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n724), .B2(new_n725), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n729), .A2(new_n727), .ZN(new_n738));
  INV_X1    g313(.A(new_n695), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n608), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n675), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT23), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G171), .B2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT90), .Z(new_n750));
  OAI211_X1 g325(.A(new_n741), .B(new_n746), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n695), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n695), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT29), .B(G2090), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n675), .A2(G21), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G286), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n692), .B1(new_n760), .B2(G28), .ZN(new_n762));
  NOR2_X1   g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  AND2_X1   g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n759), .B1(new_n761), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n695), .A2(G27), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n695), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT91), .B(G2078), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n757), .B2(new_n758), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n755), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n739), .A2(G26), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT28), .Z(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(G116), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n487), .B2(G128), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n494), .A2(G140), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n777), .A2(KEYINPUT87), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(KEYINPUT87), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n773), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2067), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n692), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  AOI22_X1  g362(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n462), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n494), .A2(G139), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n494), .A2(KEYINPUT88), .A3(G139), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n785), .B1(new_n794), .B2(new_n692), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G2072), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT89), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(G2072), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n771), .A2(new_n784), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n675), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n592), .B2(new_n675), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n750), .A2(new_n747), .B1(G1348), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G1348), .B2(new_n801), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n751), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n712), .B(new_n804), .C1(new_n710), .C2(new_n708), .ZN(G150));
  XOR2_X1   g380(.A(G150), .B(KEYINPUT93), .Z(G311));
  NAND2_X1  g381(.A1(new_n592), .A2(G559), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n534), .A2(G55), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n526), .A2(G93), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n514), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n546), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n546), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n809), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n820), .A2(new_n821), .A3(G860), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n815), .A2(G860), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  NAND2_X1  g400(.A1(new_n510), .A2(new_n507), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n502), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT96), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n779), .B2(new_n780), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n777), .A2(new_n778), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT87), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n777), .A2(KEYINPUT87), .A3(new_n778), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n830), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n721), .ZN(new_n839));
  INV_X1    g414(.A(new_n794), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n832), .A2(new_n837), .A3(new_n722), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n839), .A2(KEYINPUT98), .A3(new_n840), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n832), .A2(new_n837), .A3(new_n722), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n722), .B1(new_n832), .B2(new_n837), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n794), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT97), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT97), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n494), .A2(G142), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n487), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n462), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n701), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n849), .B(KEYINPUT97), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n846), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n614), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n852), .A2(new_n859), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n861), .A3(new_n846), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n613), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n608), .B(G160), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G162), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n864), .A2(new_n872), .A3(new_n867), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT40), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n860), .A2(new_n863), .A3(new_n614), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n613), .B1(new_n865), .B2(new_n866), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  AND4_X1   g453(.A1(KEYINPUT40), .A2(new_n877), .A3(new_n878), .A4(new_n873), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(new_n879), .ZN(G395));
  XNOR2_X1  g455(.A(new_n582), .B(G305), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n565), .B(G166), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n818), .B(new_n599), .ZN(new_n886));
  INV_X1    g461(.A(G299), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n591), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(KEYINPUT41), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n885), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n815), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n898), .ZN(G295));
  OAI21_X1  g474(.A(new_n897), .B1(G868), .B2(new_n898), .ZN(G331));
  XNOR2_X1  g475(.A(G168), .B(G301), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n818), .B(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n888), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n883), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(G37), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n904), .B(new_n883), .C1(new_n890), .C2(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT102), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n903), .A2(new_n909), .A3(new_n883), .A4(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(KEYINPUT44), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(G397));
  XOR2_X1   g495(.A(KEYINPUT103), .B(G1384), .Z(new_n921));
  AND2_X1   g496(.A1(new_n830), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT45), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n467), .A2(G40), .A3(new_n470), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n479), .B1(new_n478), .B2(G2105), .ZN(new_n925));
  AOI211_X1 g500(.A(KEYINPUT66), .B(new_n462), .C1(new_n477), .C2(new_n472), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n476), .A2(new_n480), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n924), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n781), .B(G2067), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n721), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n701), .B(new_n703), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g517(.A1(G290), .A2(G1986), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n933), .C1(new_n942), .C2(new_n943), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(G303), .A2(G8), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT106), .B(G1971), .ZN(new_n949));
  OAI21_X1  g524(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n474), .A2(new_n500), .B1(new_n951), .B2(new_n498), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n826), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(KEYINPUT45), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n922), .B2(KEYINPUT45), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n949), .B1(new_n955), .B2(new_n932), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n930), .B1(new_n929), .B2(new_n924), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n467), .A2(G40), .A3(new_n470), .ZN(new_n961));
  AOI211_X1 g536(.A(KEYINPUT104), .B(new_n961), .C1(new_n476), .C2(new_n480), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  INV_X1    g540(.A(new_n507), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n506), .B1(new_n474), .B2(new_n504), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n829), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n952), .A2(KEYINPUT96), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n964), .B(new_n965), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT107), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n830), .A2(new_n972), .A3(new_n964), .A4(new_n965), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n963), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2090), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n958), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n932), .A2(new_n959), .A3(new_n971), .A4(new_n973), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n978), .A2(KEYINPUT108), .A3(G2090), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT109), .B(new_n957), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G8), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT108), .B1(new_n978), .B2(G2090), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n971), .A2(new_n973), .ZN(new_n983));
  INV_X1    g558(.A(new_n959), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n928), .B2(new_n931), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n983), .A2(new_n985), .A3(new_n958), .A4(new_n976), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n956), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT109), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n948), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n987), .B2(KEYINPUT109), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n957), .B1(new_n977), .B2(new_n979), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n948), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n573), .A2(new_n997), .A3(new_n665), .A4(new_n574), .ZN(new_n998));
  INV_X1    g573(.A(new_n569), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT75), .B1(new_n571), .B2(new_n514), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n574), .A2(new_n665), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT111), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n572), .B1(KEYINPUT112), .B2(new_n569), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n569), .A2(KEYINPUT112), .ZN(new_n1005));
  OAI21_X1  g580(.A(G1981), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n830), .A2(new_n965), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n990), .B1(new_n932), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1003), .B(new_n1006), .C1(KEYINPUT113), .C2(KEYINPUT49), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n677), .A2(G1976), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT110), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1024), .A3(new_n1018), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1019), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1010), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n960), .B2(new_n962), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT114), .B1(new_n953), .B2(KEYINPUT45), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  NOR4_X1   g606(.A1(G164), .A2(new_n1031), .A3(new_n1027), .A4(G1384), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n758), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1035));
  INV_X1    g610(.A(G2084), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n983), .A2(new_n1036), .A3(new_n985), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n758), .C1(new_n1029), .C2(new_n1033), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n989), .A2(new_n996), .A3(new_n1026), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n991), .A2(new_n994), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(new_n948), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n996), .A4(new_n1026), .ZN(new_n1048));
  INV_X1    g623(.A(new_n932), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n953), .A2(new_n964), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1011), .B2(new_n964), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1049), .A2(new_n1051), .A3(G2090), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1052), .B2(new_n956), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n948), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1040), .A2(G8), .A3(G168), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n996), .A2(new_n1026), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1044), .A2(new_n1048), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n996), .A2(new_n1026), .A3(new_n1054), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n975), .A2(KEYINPUT119), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n978), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1064), .A3(new_n747), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n955), .A2(new_n1066), .A3(new_n932), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n932), .B(new_n1028), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1065), .B(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G171), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1061), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1039), .A2(new_n1037), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1038), .B1(new_n1070), .B2(new_n758), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT124), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1035), .A2(new_n1078), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(G168), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n990), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1040), .A2(G8), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G286), .A2(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT62), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1080), .A2(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1089), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1074), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1060), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1026), .A2(new_n995), .A3(new_n994), .A4(new_n991), .ZN(new_n1097));
  AOI211_X1 g672(.A(G1976), .B(G288), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1003), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1012), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(G1996), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n955), .A2(new_n932), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n932), .A2(new_n1011), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  AOI22_X1  g681(.A1(new_n1103), .A2(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n955), .A2(KEYINPUT121), .A3(new_n932), .A4(new_n1102), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n546), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT59), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n547), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1111), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1110), .A2(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1348), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1062), .A2(new_n1064), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G2067), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n932), .A2(new_n1125), .A3(new_n1011), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n592), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n555), .B2(new_n559), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT117), .B(G1956), .Z(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(G2072), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n955), .A2(new_n932), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT61), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1132), .B2(new_n1130), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1139), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1128), .A2(new_n1129), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1112), .A2(new_n1119), .A3(new_n1110), .A4(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n591), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1122), .A2(new_n1147), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n592), .A3(new_n1139), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1144), .A3(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(G301), .B(KEYINPUT54), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1066), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n478), .B2(G2105), .ZN(new_n1158));
  INV_X1    g733(.A(new_n471), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(KEYINPUT125), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1160), .B(new_n923), .C1(KEYINPUT125), .C2(new_n1159), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT45), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1155), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1155), .A2(new_n1072), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1092), .B2(new_n1089), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1061), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1101), .B1(new_n1154), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n946), .B1(new_n1096), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n937), .A2(new_n933), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n701), .A2(new_n703), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1169), .A2(new_n1170), .B1(new_n1125), .B2(new_n781), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n933), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n935), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT46), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n722), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n933), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n933), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT48), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n939), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1175), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT127), .B1(new_n1168), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n946), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1101), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1153), .A2(new_n1144), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1152), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1165), .A2(new_n1061), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1060), .A2(new_n1095), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1186), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1184), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1185), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g772(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n672), .A2(new_n1199), .A3(new_n673), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n913), .B2(new_n915), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n871), .A2(new_n873), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1202), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


