//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n914, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT1), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(G127gat), .A2(G134gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G127gat), .A2(G134gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G113gat), .B(G120gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n212), .B(KEYINPUT68), .C1(new_n213), .C2(KEYINPUT1), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n204), .A2(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT69), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(new_n208), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(G155gat), .B2(G162gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G148gat), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G141gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G155gat), .B(G162gat), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT2), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n229), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n229), .A2(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n215), .A2(new_n240), .A3(new_n221), .A4(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n208), .A2(new_n220), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n204), .A2(new_n206), .A3(new_n218), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n217), .A2(new_n254), .B1(new_n209), .B2(new_n214), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n255), .A2(KEYINPUT79), .A3(new_n248), .A4(new_n240), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n215), .A2(new_n240), .A3(new_n221), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n246), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n215), .A2(new_n240), .A3(new_n221), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n240), .B1(new_n221), .B2(new_n215), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT80), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n222), .A2(new_n243), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n257), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT80), .A3(new_n261), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(KEYINPUT5), .A3(new_n266), .A4(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n271));
  INV_X1    g070(.A(new_n258), .ZN(new_n272));
  INV_X1    g071(.A(new_n249), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n245), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G57gat), .B(G85gat), .Z(new_n276));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT40), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n258), .A2(new_n249), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n246), .B1(new_n284), .B2(new_n245), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT39), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT39), .B1(new_n268), .B2(new_n261), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n282), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n283), .B2(new_n289), .ZN(new_n291));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT22), .ZN(new_n293));
  INV_X1    g092(.A(G211gat), .ZN(new_n294));
  INV_X1    g093(.A(G218gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n292), .A3(new_n296), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT65), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT25), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  AOI211_X1 g124(.A(KEYINPUT65), .B(new_n325), .C1(new_n313), .C2(new_n321), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n314), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n310), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n307), .B1(new_n329), .B2(KEYINPUT26), .ZN(new_n330));
  NOR2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT26), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n328), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G183gat), .ZN(new_n336));
  AOI21_X1  g135(.A(G190gat), .B1(new_n336), .B2(KEYINPUT27), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n338), .A3(G183gat), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT28), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT27), .B(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G190gat), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n334), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n327), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT76), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n312), .ZN(new_n351));
  NOR3_X1   g150(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n323), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n325), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT25), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n345), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n348), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT27), .B1(new_n318), .B2(KEYINPUT66), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n339), .A3(new_n319), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n369));
  INV_X1    g168(.A(new_n333), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n350), .B1(new_n331), .B2(new_n332), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n314), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT67), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT67), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n334), .B(new_n374), .C1(new_n340), .C2(new_n344), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n327), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n327), .A3(KEYINPUT74), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n347), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n306), .B1(new_n366), .B2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n348), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n379), .B2(new_n380), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n361), .A2(new_n347), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n305), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT77), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n382), .A2(new_n388), .A3(new_n395), .A4(new_n392), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n388), .ZN(new_n398));
  INV_X1    g197(.A(new_n392), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT30), .B(new_n392), .C1(new_n382), .C2(new_n388), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n394), .B(new_n396), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT88), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n394), .A2(new_n396), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n363), .A2(new_n364), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT76), .B(new_n348), .C1(new_n361), .C2(new_n362), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n380), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT74), .B1(new_n376), .B2(new_n327), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n348), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n305), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n384), .B1(new_n409), .B2(new_n410), .ZN(new_n413));
  INV_X1    g212(.A(new_n387), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n306), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n399), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT30), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n392), .B1(new_n382), .B2(new_n388), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n397), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n291), .B1(new_n403), .B2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT85), .B(G78gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G22gat), .B(G50gat), .Z(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n383), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n242), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n305), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT87), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n433), .A3(new_n305), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n303), .A2(new_n362), .A3(new_n243), .A4(new_n304), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n244), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT86), .ZN(new_n438));
  INV_X1    g237(.A(G228gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n437), .A2(KEYINPUT86), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n438), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G106gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n431), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n300), .A2(new_n302), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n429), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n240), .B1(new_n447), .B2(new_n241), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n445), .A2(new_n448), .B1(new_n439), .B2(new_n440), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n443), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n428), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n450), .A3(new_n427), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n280), .B1(new_n270), .B2(new_n274), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT90), .B1(new_n457), .B2(KEYINPUT6), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(KEYINPUT6), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT5), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n247), .A2(new_n259), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n280), .B(new_n274), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n465), .B2(KEYINPUT90), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n412), .B2(new_n415), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n382), .A2(KEYINPUT37), .A3(new_n388), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n392), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n418), .B1(new_n470), .B2(KEYINPUT38), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n408), .A2(new_n305), .A3(new_n411), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n413), .A2(new_n306), .A3(new_n414), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT37), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n468), .A2(new_n472), .A3(new_n392), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n399), .B1(new_n398), .B2(new_n467), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n472), .A4(new_n475), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n466), .A2(new_n471), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n422), .A2(new_n456), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n462), .A2(new_n484), .A3(new_n463), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n282), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n459), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(KEYINPUT83), .A3(new_n420), .A4(new_n405), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n489));
  INV_X1    g288(.A(new_n459), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n457), .B1(new_n464), .B2(KEYINPUT82), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n485), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n489), .B1(new_n492), .B2(new_n402), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n456), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n377), .A2(new_n222), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n376), .A2(new_n327), .A3(new_n255), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(KEYINPUT64), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT33), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT70), .B(G15gat), .ZN(new_n510));
  INV_X1    g309(.A(G43gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G71gat), .B(G99gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n507), .A2(KEYINPUT32), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n509), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n506), .A2(KEYINPUT34), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n502), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n522));
  AOI22_X1  g321(.A1(KEYINPUT71), .A2(new_n521), .B1(new_n522), .B2(KEYINPUT34), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n516), .A2(new_n524), .A3(new_n523), .A4(new_n518), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n499), .B(new_n500), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(new_n525), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(new_n527), .A3(new_n497), .A4(new_n498), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n482), .A2(new_n496), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n456), .A2(new_n530), .A3(new_n527), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n488), .A2(new_n493), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n403), .A2(new_n421), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT35), .ZN(new_n539));
  INV_X1    g338(.A(new_n466), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n535), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(G1gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT93), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n544), .A2(G1gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(KEYINPUT93), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(G8gat), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n546), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G8gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(G57gat), .A2(G64gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G57gat), .A2(G64gat), .ZN(new_n556));
  AND2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT100), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(new_n557), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n554), .B1(KEYINPUT21), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT101), .ZN(new_n565));
  AND2_X1   g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n563), .A2(KEYINPUT21), .ZN(new_n569));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  OAI21_X1  g376(.A(new_n572), .B1(new_n567), .B2(new_n568), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n574), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT103), .ZN(new_n583));
  XOR2_X1   g382(.A(G43gat), .B(G50gat), .Z(new_n584));
  XOR2_X1   g383(.A(KEYINPUT91), .B(G36gat), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G29gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT14), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(G29gat), .B2(G36gat), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n587), .A2(G29gat), .A3(G36gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT15), .ZN(new_n590));
  INV_X1    g389(.A(G50gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(G43gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n592), .B2(KEYINPUT92), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n584), .A2(new_n594), .B1(new_n595), .B2(new_n590), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n594), .A2(new_n584), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT17), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT7), .ZN(new_n601));
  INV_X1    g400(.A(G99gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT8), .B1(new_n602), .B2(new_n444), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n603), .C1(G85gat), .C2(G92gat), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n598), .A2(KEYINPUT17), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n598), .A2(new_n606), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(KEYINPUT41), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n612), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n583), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n619), .A2(new_n620), .A3(new_n583), .ZN(new_n623));
  OAI22_X1  g422(.A1(new_n622), .A2(new_n623), .B1(new_n614), .B2(new_n613), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n613), .A2(new_n614), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n621), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n581), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n598), .B(new_n554), .Z(new_n631));
  XOR2_X1   g430(.A(KEYINPUT98), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(G229gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT99), .Z(new_n636));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n554), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n599), .A3(new_n607), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n598), .B1(new_n553), .B2(new_n551), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n641), .A2(new_n643), .A3(KEYINPUT18), .A4(new_n633), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n633), .A3(new_n643), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n649));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650));
  INV_X1    g449(.A(G197gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT11), .B(G169gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n645), .B(new_n648), .C1(new_n649), .C2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n636), .A2(new_n649), .A3(new_n644), .ZN(new_n657));
  INV_X1    g456(.A(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n644), .ZN(new_n659));
  INV_X1    g458(.A(new_n648), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n657), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n606), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n563), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n606), .A2(new_n562), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT104), .A4(new_n666), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n663), .A2(KEYINPUT10), .A3(new_n563), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n664), .A2(new_n665), .ZN(new_n675));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n677), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n682), .A2(KEYINPUT105), .A3(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n662), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n630), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n543), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n492), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(new_n538), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT16), .B(G8gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT42), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(G8gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1325gat));
  OAI21_X1  g502(.A(G15gat), .B1(new_n692), .B2(new_n533), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n526), .A2(new_n528), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n692), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT107), .Z(G1326gat));
  NOR2_X1   g508(.A1(new_n692), .A2(new_n456), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(new_n581), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n690), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n543), .A2(new_n628), .A3(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n487), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT45), .Z(new_n717));
  AND2_X1   g516(.A1(new_n481), .A2(new_n456), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n532), .B1(new_n718), .B2(new_n422), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n719), .A2(new_n496), .B1(new_n537), .B2(new_n541), .ZN(new_n720));
  INV_X1    g519(.A(new_n628), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT44), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n543), .A2(new_n723), .A3(new_n628), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n714), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n487), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n727), .ZN(G1328gat));
  NOR3_X1   g527(.A1(new_n715), .A2(new_n538), .A3(new_n585), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n585), .B1(new_n726), .B2(new_n538), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1329gat));
  OAI21_X1  g531(.A(G43gat), .B1(new_n726), .B2(new_n533), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n705), .A2(new_n511), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n715), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g535(.A1(new_n456), .A2(new_n591), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n723), .B1(new_n543), .B2(new_n628), .ZN(new_n738));
  AOI211_X1 g537(.A(KEYINPUT44), .B(new_n721), .C1(new_n534), .C2(new_n542), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n714), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n591), .B1(new_n715), .B2(new_n456), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n741), .A4(new_n742), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n742), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT109), .B1(new_n748), .B2(KEYINPUT48), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n750), .B(new_n741), .C1(new_n740), .C2(new_n742), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n745), .A2(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n743), .A2(new_n744), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n746), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n755), .B(new_n756), .C1(new_n749), .C2(new_n751), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(G1331gat));
  NOR3_X1   g557(.A1(new_n630), .A2(new_n662), .A3(new_n689), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n543), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n492), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G57gat), .ZN(G1332gat));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n764));
  INV_X1    g563(.A(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n696), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n765), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n760), .B2(new_n533), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n706), .A2(G71gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n760), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n761), .A2(new_n495), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  INV_X1    g576(.A(new_n689), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n713), .A2(new_n662), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n725), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(G85gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n487), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n543), .A2(new_n628), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n785), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n492), .A3(new_n778), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n782), .B1(new_n790), .B2(new_n781), .ZN(G1336gat));
  NOR2_X1   g590(.A1(new_n780), .A2(new_n538), .ZN(new_n792));
  INV_X1    g591(.A(G92gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n783), .B(new_n795), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n538), .A2(G92gat), .A3(new_n689), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n789), .A2(new_n778), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(G92gat), .A3(new_n538), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n792), .B2(new_n793), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n798), .A2(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n780), .B2(new_n533), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n705), .A2(new_n602), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n800), .B2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n689), .A2(G106gat), .A3(new_n456), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n780), .A2(new_n456), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n444), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n444), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n807), .B(KEYINPUT115), .Z(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n796), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n814), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g614(.A(new_n662), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n629), .A2(new_n816), .A3(new_n689), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n648), .A2(new_n636), .A3(new_n644), .A4(new_n655), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n633), .B1(new_n641), .B2(new_n643), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n631), .A2(new_n634), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n654), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n627), .B(new_n624), .C1(new_n689), .C2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n681), .B1(new_n674), .B2(KEYINPUT54), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n669), .A2(new_n676), .A3(new_n670), .A4(new_n671), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n826), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n824), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n831), .A3(new_n684), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n656), .B2(new_n661), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n581), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(KEYINPUT116), .B2(new_n822), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n721), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n817), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n696), .A2(new_n487), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT117), .B(new_n817), .C1(new_n834), .C2(new_n837), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n840), .A2(new_n535), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n816), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n662), .A2(new_n205), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT118), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n843), .B2(new_n846), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n843), .A2(new_n689), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n203), .ZN(G1341gat));
  NOR2_X1   g648(.A1(new_n843), .A2(new_n581), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g650(.A1(new_n843), .A2(new_n721), .ZN(new_n852));
  INV_X1    g651(.A(G134gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n857), .A3(new_n853), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n858), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n855), .A2(new_n863), .A3(new_n856), .A4(new_n858), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n843), .B2(new_n721), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n860), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(G1343gat));
  NAND3_X1  g665(.A1(new_n840), .A2(new_n495), .A3(new_n842), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n533), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n230), .A3(new_n662), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n838), .A2(KEYINPUT57), .A3(new_n495), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  XOR2_X1   g671(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n816), .A3(new_n868), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n870), .B1(new_n876), .B2(new_n230), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n232), .A3(new_n778), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT122), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n875), .A2(new_n689), .A3(new_n868), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n232), .A2(KEYINPUT59), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n868), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n867), .A2(new_n874), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n778), .B(new_n886), .C1(new_n887), .C2(new_n872), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(KEYINPUT123), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n840), .A2(new_n495), .A3(new_n842), .A4(new_n873), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n838), .A2(new_n495), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n892), .B2(new_n893), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n778), .B(new_n886), .C1(new_n895), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n891), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n880), .B1(new_n890), .B2(new_n901), .ZN(G1345gat));
  AOI21_X1  g701(.A(G155gat), .B1(new_n869), .B2(new_n713), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n875), .A2(new_n868), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n581), .A2(new_n236), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n869), .A2(new_n237), .A3(new_n628), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n875), .A2(new_n721), .A3(new_n868), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n237), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n538), .A2(new_n492), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n840), .A2(new_n535), .A3(new_n842), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n816), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(new_n309), .ZN(G1348gat));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n689), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(new_n310), .ZN(G1349gat));
  OAI21_X1  g714(.A(new_n318), .B1(new_n911), .B2(new_n581), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n911), .A2(new_n581), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n341), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT60), .Z(G1350gat));
  NOR2_X1   g718(.A1(new_n911), .A2(new_n721), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n319), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT61), .B(G190gat), .Z(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n920), .B2(new_n923), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n532), .A2(new_n538), .A3(new_n492), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n840), .A2(new_n495), .A3(new_n842), .A4(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n651), .B(new_n662), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n895), .A2(new_n899), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n925), .B(KEYINPUT126), .Z(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT127), .Z(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n662), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n930), .B1(new_n935), .B2(new_n651), .ZN(G1352gat));
  NAND3_X1  g735(.A1(new_n931), .A2(new_n778), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G204gat), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n689), .A2(G204gat), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT62), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n926), .A2(KEYINPUT62), .A3(new_n939), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(G1353gat));
  OAI211_X1 g741(.A(new_n294), .B(new_n713), .C1(new_n928), .C2(new_n929), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n713), .B(new_n932), .C1(new_n895), .C2(new_n899), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  AND2_X1   g746(.A1(new_n931), .A2(new_n933), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n721), .A2(new_n295), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n628), .B1(new_n928), .B2(new_n929), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n948), .A2(new_n949), .B1(new_n295), .B2(new_n950), .ZN(G1355gat));
endmodule


