//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1184, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND3_X1  g0006(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(new_n203), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n208), .A2(new_n210), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g0015(.A1(G87), .A2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT67), .B(G244), .Z(new_n221));
  AOI211_X1 g0021(.A(new_n216), .B(new_n220), .C1(new_n221), .C2(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT66), .B(G238), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n203), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n215), .B(new_n229), .C1(new_n211), .C2(new_n214), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n223), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  INV_X1    g0033(.A(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G107), .ZN(new_n244));
  INV_X1    g0044(.A(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G351));
  XOR2_X1   g0047(.A(KEYINPUT8), .B(G58), .Z(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n204), .A2(G20), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n248), .A2(new_n250), .B1(new_n251), .B2(KEYINPUT72), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n252), .B1(KEYINPUT72), .B2(new_n251), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n256), .A2(new_n259), .B1(new_n201), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n261), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n259), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G50), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G223), .A3(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(G222), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G77), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n270), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT70), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n258), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n270), .A2(new_n272), .A3(KEYINPUT70), .A4(new_n276), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n260), .B(G274), .C1(G41), .C2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT68), .B(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(new_n283), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT71), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n282), .A2(new_n294), .A3(new_n283), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n268), .B1(new_n296), .B2(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(G179), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n269), .A2(G232), .A3(new_n271), .ZN(new_n300));
  INV_X1    g0100(.A(G107), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n269), .A2(G1698), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n300), .B1(new_n301), .B2(new_n269), .C1(new_n302), .C2(new_n224), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n280), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n289), .A2(new_n221), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n283), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(G179), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n263), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT73), .ZN(new_n312));
  INV_X1    g0112(.A(new_n266), .ZN(new_n313));
  INV_X1    g0113(.A(new_n248), .ZN(new_n314));
  INV_X1    g0114(.A(G20), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n314), .A2(new_n255), .B1(new_n315), .B2(new_n310), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n250), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n259), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n312), .B1(new_n310), .B2(new_n313), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n307), .A2(new_n309), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n306), .B2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n306), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n299), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n248), .A2(new_n261), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT76), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n263), .A2(new_n259), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n314), .A2(new_n263), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT75), .B1(new_n202), .B2(new_n203), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G58), .A3(G68), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n337), .A3(new_n209), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(G159), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n255), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n315), .ZN(new_n342));
  OR2_X1    g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT74), .B1(new_n273), .B2(new_n274), .ZN(new_n347));
  AOI21_X1  g0147(.A(G20), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n342), .B1(new_n348), .B2(KEYINPUT7), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n341), .B1(new_n349), .B2(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n320), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n275), .B2(new_n315), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n203), .B1(new_n354), .B2(new_n342), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n352), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n334), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n285), .A2(G232), .A3(new_n286), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n358), .A2(KEYINPUT78), .A3(new_n283), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT78), .B1(new_n358), .B2(new_n283), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(G226), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n362));
  OAI211_X1 g0162(.A(G223), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT77), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n361), .B1(new_n369), .B2(new_n280), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n285), .B1(new_n367), .B2(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n358), .A2(new_n283), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n308), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n328), .B1(new_n357), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n338), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n269), .A2(new_n379), .A3(G20), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT74), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n315), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT16), .B(new_n378), .C1(new_n384), .C2(new_n203), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n356), .A3(new_n259), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n332), .A2(new_n333), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n369), .A2(new_n280), .ZN(new_n389));
  INV_X1    g0189(.A(new_n374), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n308), .B1(new_n370), .B2(new_n371), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n392), .A3(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n377), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G200), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n391), .A2(new_n395), .B1(new_n370), .B2(new_n324), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT17), .B1(new_n388), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n370), .A2(new_n324), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n395), .B1(new_n373), .B2(new_n374), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n357), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n394), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n296), .A2(G190), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n293), .A2(G200), .A3(new_n295), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n268), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n407), .A2(new_n409), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT10), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n406), .A4(new_n405), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n404), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n289), .A2(G238), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n269), .A2(G232), .A3(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n269), .A2(new_n271), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n418), .C1(new_n419), .C2(new_n234), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n280), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n283), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT14), .B1(new_n425), .B2(new_n308), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(G179), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(G169), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n250), .A2(G77), .B1(new_n254), .B2(G50), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n315), .B2(G68), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n203), .B2(new_n313), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n263), .A2(new_n203), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT12), .Z(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT11), .B1(new_n432), .B2(new_n259), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n425), .B2(new_n395), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n423), .A2(new_n424), .A3(new_n324), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n327), .A2(new_n415), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT79), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n448));
  OAI211_X1 g0248(.A(G250), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G294), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n280), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n260), .A2(G45), .ZN(new_n453));
  OR2_X1    g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n280), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G264), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(G274), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n452), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT84), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n460), .A2(new_n461), .A3(new_n395), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n460), .B2(new_n395), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n460), .A2(G190), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n315), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n269), .A2(new_n469), .A3(new_n315), .A4(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n249), .A2(new_n245), .A3(G20), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n315), .A2(G107), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT23), .ZN(new_n475));
  AND4_X1   g0275(.A1(new_n466), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n468), .B2(new_n470), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n466), .B1(new_n477), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n259), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n260), .A2(G33), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n331), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n301), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n263), .A2(new_n301), .ZN(new_n484));
  XOR2_X1   g0284(.A(new_n484), .B(KEYINPUT25), .Z(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n465), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n452), .A2(new_n458), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n371), .A3(new_n459), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n460), .A2(new_n308), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n477), .A2(new_n466), .A3(new_n475), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n482), .B1(new_n495), .B2(new_n259), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n491), .B1(new_n496), .B2(new_n485), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT85), .B1(new_n487), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n460), .A2(new_n395), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT84), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n460), .A2(new_n461), .A3(new_n395), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n496), .B(new_n485), .C1(new_n502), .C2(new_n464), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G244), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n269), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n280), .ZN(new_n515));
  INV_X1    g0315(.A(G45), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(G1), .ZN(new_n517));
  INV_X1    g0317(.A(new_n455), .ZN(new_n518));
  NOR2_X1   g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n285), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n459), .B1(new_n521), .B2(new_n219), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n515), .A2(new_n523), .A3(new_n371), .ZN(new_n524));
  AOI21_X1  g0324(.A(G169), .B1(new_n515), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT81), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n265), .A2(G13), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(G97), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n380), .B2(new_n353), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n301), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n218), .A2(new_n301), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n533), .B2(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n254), .A2(G77), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n528), .B1(new_n537), .B2(new_n259), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n218), .B2(new_n481), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n515), .A2(new_n523), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G179), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n526), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n269), .A2(G244), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n269), .A2(G238), .A3(new_n271), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(new_n545), .C1(new_n249), .C2(new_n245), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n280), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n517), .A2(G274), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n285), .A2(G250), .A3(new_n453), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n547), .A2(new_n371), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n315), .B1(new_n418), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n532), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n315), .A2(G33), .A3(G97), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n552), .A2(new_n554), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n269), .A2(new_n315), .A3(G68), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n320), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n318), .A2(new_n527), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n317), .B(KEYINPUT82), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n527), .A2(new_n320), .A3(new_n480), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n548), .ZN(new_n565));
  INV_X1    g0365(.A(new_n549), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n546), .C2(new_n280), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n550), .B(new_n564), .C1(new_n567), .C2(G169), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n547), .A2(G190), .A3(new_n548), .A4(new_n549), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n481), .A2(new_n553), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n570), .A2(new_n558), .A3(new_n559), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n571), .C1(new_n567), .C2(new_n395), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT80), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n541), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n522), .B1(new_n280), .B2(new_n514), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(G200), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n481), .A2(new_n218), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n528), .B(new_n579), .C1(new_n537), .C2(new_n259), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(G190), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n543), .A2(new_n573), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n562), .A2(G116), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n512), .B(new_n315), .C1(G33), .C2(new_n218), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n259), .C1(new_n315), .C2(G116), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  OAI221_X1 g0390(.A(new_n585), .B1(G116), .B2(new_n527), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n269), .A2(G264), .A3(G1698), .ZN(new_n592));
  INV_X1    g0392(.A(G303), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n592), .B1(new_n593), .B2(new_n269), .C1(new_n419), .C2(new_n219), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n280), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n457), .A2(G270), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n459), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n597), .A3(G169), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(new_n371), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n591), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n591), .A2(new_n597), .A3(KEYINPUT21), .A4(G169), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(G200), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n324), .B2(new_n597), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n591), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n543), .A2(new_n573), .A3(new_n582), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT83), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n507), .A2(new_n584), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n447), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT86), .ZN(G372));
  INV_X1    g0413(.A(new_n572), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n550), .A2(new_n564), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT87), .B1(new_n567), .B2(G169), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n308), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n614), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n526), .A2(KEYINPUT88), .A3(new_n542), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT88), .B1(new_n526), .B2(new_n542), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n539), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n543), .B(new_n582), .C1(new_n604), .C2(new_n497), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n503), .ZN(new_n626));
  OAI22_X1  g0426(.A1(new_n624), .A2(KEYINPUT26), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n620), .A2(new_n615), .ZN(new_n628));
  INV_X1    g0428(.A(new_n573), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n543), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n446), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n299), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT89), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT89), .B1(new_n411), .B2(new_n414), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n440), .A2(new_n322), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n444), .A2(new_n403), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n394), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n635), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n634), .A2(new_n642), .ZN(G369));
  XNOR2_X1  g0443(.A(new_n608), .B(KEYINPUT90), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n262), .A2(G20), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n260), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n591), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n604), .B2(new_n652), .ZN(new_n654));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n486), .A2(new_n651), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n507), .A2(new_n657), .B1(new_n497), .B2(new_n651), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n651), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n604), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n498), .B2(new_n506), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n497), .B2(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n213), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n554), .A2(G116), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n210), .B2(new_n668), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n633), .A2(new_n661), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(KEYINPUT29), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n567), .A2(new_n488), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n601), .A2(new_n675), .A3(new_n576), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n567), .B(KEYINPUT91), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n597), .A2(new_n371), .A3(new_n460), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n541), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n601), .A2(new_n675), .A3(KEYINPUT30), .A4(new_n576), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n678), .A2(new_n681), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n651), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n611), .B2(KEYINPUT31), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n655), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n625), .A2(new_n626), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n628), .A2(KEYINPUT93), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n628), .A2(KEYINPUT93), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n630), .B2(new_n631), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n695), .B1(new_n701), .B2(new_n661), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n674), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n672), .B1(new_n703), .B2(G1), .ZN(G364));
  AOI21_X1  g0504(.A(new_n260), .B1(new_n645), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n667), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n654), .A2(new_n655), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n656), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n262), .A2(new_n249), .A3(KEYINPUT95), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT95), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G13), .B2(G33), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n654), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n242), .A2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  INV_X1    g0519(.A(new_n210), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n718), .A2(new_n719), .B1(new_n516), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n381), .A2(new_n382), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n666), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n721), .B(new_n723), .C1(new_n719), .C2(new_n718), .ZN(new_n724));
  INV_X1    g0524(.A(G355), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n269), .A2(new_n213), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n724), .B1(G116), .B2(new_n213), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n258), .B1(G20), .B2(new_n308), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n716), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n315), .A2(new_n371), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n269), .B1(new_n733), .B2(G326), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n324), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G317), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT33), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(KEYINPUT33), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n315), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n395), .A2(G179), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n734), .B(new_n740), .C1(new_n741), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n315), .A2(new_n324), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n371), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G322), .A2(new_n749), .B1(new_n752), .B2(G329), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n746), .A2(new_n743), .ZN(new_n754));
  INV_X1    g0554(.A(G311), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n742), .A2(new_n747), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n753), .B1(new_n593), .B2(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n315), .B1(new_n750), .B2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n745), .B(new_n757), .C1(G294), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n754), .ZN(new_n761));
  INV_X1    g0561(.A(new_n756), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G87), .A2(new_n761), .B1(new_n762), .B2(G77), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n763), .B1(new_n202), .B2(new_n748), .C1(new_n301), .C2(new_n744), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT96), .B(G159), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n752), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT32), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n735), .A2(new_n203), .B1(new_n758), .B2(new_n218), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n269), .B1(new_n732), .B2(new_n201), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n764), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n728), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n717), .A2(new_n707), .A3(new_n730), .A4(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n710), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(G396));
  NOR2_X1   g0574(.A1(new_n322), .A2(new_n651), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n321), .A2(new_n651), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n325), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(new_n777), .B2(new_n322), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n673), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n661), .C1(new_n627), .C2(new_n632), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(new_n694), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n708), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n735), .A2(new_n741), .B1(new_n732), .B2(new_n593), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G97), .B2(new_n759), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n749), .A2(G294), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n754), .A2(new_n301), .B1(new_n751), .B2(new_n755), .ZN(new_n788));
  INV_X1    g0588(.A(new_n744), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G87), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n269), .B1(new_n762), .B2(G116), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n787), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n733), .A2(G137), .B1(new_n762), .B2(new_n765), .ZN(new_n793));
  INV_X1    g0593(.A(G143), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n794), .B2(new_n748), .C1(new_n253), .C2(new_n735), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT34), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n754), .A2(new_n201), .B1(new_n744), .B2(new_n203), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT97), .ZN(new_n800));
  INV_X1    g0600(.A(new_n722), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G58), .B2(new_n759), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n797), .A2(new_n798), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n752), .A2(G132), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n792), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n714), .A2(new_n728), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n805), .A2(new_n728), .B1(new_n310), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n707), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT98), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n715), .B2(new_n778), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n784), .A2(new_n810), .ZN(G384));
  NAND2_X1  g0611(.A1(new_n439), .A2(new_n651), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n440), .A2(new_n444), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n439), .B(new_n651), .C1(new_n430), .C2(new_n443), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n690), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n778), .B(new_n815), .C1(new_n687), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT101), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n649), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n388), .B1(new_n392), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n357), .A2(new_n401), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT37), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n350), .A2(KEYINPUT16), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n334), .B1(new_n824), .B2(new_n351), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n820), .B1(new_n372), .B2(new_n375), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n822), .B(KEYINPUT37), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n649), .B1(new_n394), .B2(new_n403), .ZN(new_n829));
  INV_X1    g0629(.A(new_n825), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n823), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT99), .B1(new_n831), .B2(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  INV_X1    g0633(.A(new_n823), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT38), .A4(new_n827), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n827), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n832), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n608), .A2(new_n584), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n498), .A2(new_n506), .B1(new_n609), .B2(KEYINPUT83), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n682), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n690), .B1(new_n843), .B2(new_n686), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n844), .A2(KEYINPUT101), .A3(new_n778), .A4(new_n815), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n819), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT40), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(KEYINPUT102), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n817), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n388), .A2(new_n820), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT100), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n821), .A2(new_n822), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n854), .B1(new_n394), .B2(new_n403), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n838), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n835), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n853), .A2(KEYINPUT40), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n446), .A2(new_n844), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n863), .B(new_n864), .Z(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G330), .ZN(new_n866));
  INV_X1    g0666(.A(new_n775), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n781), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n840), .A2(new_n815), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(KEYINPUT39), .B2(new_n840), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n430), .A2(new_n439), .A3(new_n661), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n869), .B1(new_n394), .B2(new_n820), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n446), .B1(new_n702), .B2(new_n674), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n642), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n873), .B(new_n875), .Z(new_n876));
  XNOR2_X1  g0676(.A(new_n866), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n260), .B2(new_n645), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n245), .B1(new_n534), .B2(KEYINPUT35), .ZN(new_n879));
  INV_X1    g0679(.A(new_n208), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n879), .B(new_n880), .C1(KEYINPUT35), .C2(new_n534), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT36), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n720), .A2(G77), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n335), .A2(new_n337), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n883), .A2(new_n884), .B1(G50), .B2(new_n203), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(G1), .A3(new_n262), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n878), .A2(new_n882), .A3(new_n886), .ZN(G367));
  AND2_X1   g0687(.A1(new_n543), .A2(new_n582), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n580), .B2(new_n661), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n539), .B1(new_n622), .B2(new_n623), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n661), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n659), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n571), .A2(new_n661), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n628), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n621), .B2(new_n894), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n663), .A2(new_n888), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n891), .A2(new_n497), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n651), .B1(new_n901), .B2(new_n543), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n892), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n904), .B(new_n905), .Z(new_n906));
  XNOR2_X1  g0706(.A(new_n667), .B(KEYINPUT41), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n663), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n658), .A2(new_n662), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n656), .B(new_n913), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n703), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n660), .A2(KEYINPUT103), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n664), .A2(new_n891), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT45), .Z(new_n919));
  NOR2_X1   g0719(.A1(new_n664), .A2(new_n891), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT44), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n660), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n659), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n917), .B(new_n922), .C1(KEYINPUT103), .C2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n908), .B1(new_n925), .B2(new_n703), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n906), .B1(new_n926), .B2(new_n706), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n732), .A2(new_n755), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n928), .B(new_n722), .C1(G294), .C2(new_n736), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n749), .A2(G303), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n756), .A2(new_n741), .B1(new_n758), .B2(new_n301), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT105), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n744), .A2(new_n218), .B1(new_n751), .B2(new_n737), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n245), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT46), .B1(new_n754), .B2(new_n245), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n929), .A2(new_n930), .A3(new_n932), .A4(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G150), .A2(new_n749), .B1(new_n762), .B2(G50), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n202), .B2(new_n754), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT106), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n269), .B1(new_n744), .B2(new_n310), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n758), .A2(new_n203), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n732), .A2(new_n794), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(new_n736), .C2(new_n765), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n942), .B(new_n945), .C1(new_n940), .C2(new_n941), .ZN(new_n946));
  INV_X1    g0746(.A(G137), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n751), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n937), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n708), .B1(new_n950), .B2(new_n728), .ZN(new_n951));
  INV_X1    g0751(.A(new_n723), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n729), .B1(new_n213), .B2(new_n317), .C1(new_n238), .C2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n716), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n951), .B(new_n953), .C1(new_n954), .C2(new_n897), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n927), .A2(KEYINPUT107), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT107), .B1(new_n927), .B2(new_n955), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(G387));
  OR2_X1    g0760(.A1(new_n914), .A2(new_n703), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(new_n667), .A3(new_n915), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n752), .A2(G326), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n801), .B(new_n963), .C1(new_n245), .C2(new_n744), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT114), .ZN(new_n965));
  INV_X1    g0765(.A(G322), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n735), .A2(new_n755), .B1(new_n732), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT110), .Z(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n593), .B2(new_n756), .C1(new_n737), .C2(new_n748), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT48), .ZN(new_n970));
  INV_X1    g0770(.A(G294), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n969), .A2(new_n970), .B1(new_n971), .B2(new_n754), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G283), .B2(new_n759), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT111), .Z(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n970), .B2(new_n969), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT112), .B(KEYINPUT113), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT49), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n965), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n964), .A2(KEYINPUT114), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n975), .C2(new_n977), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n751), .A2(new_n253), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n761), .A2(G77), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n201), .B2(new_n748), .C1(new_n218), .C2(new_n744), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n801), .B(new_n983), .C1(G159), .C2(new_n733), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n314), .A2(new_n735), .B1(new_n203), .B2(new_n756), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT109), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n561), .A2(new_n759), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n980), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n708), .B1(new_n989), .B2(new_n728), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n235), .A2(new_n516), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n669), .B(new_n516), .C1(new_n203), .C2(new_n310), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT50), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n314), .B2(G50), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n248), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n991), .A2(new_n952), .A3(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n726), .A2(new_n669), .B1(G107), .B2(new_n213), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT108), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n729), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n658), .A2(new_n716), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n990), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n914), .A2(new_n706), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n962), .A2(new_n1002), .A3(new_n1003), .ZN(G393));
  NAND3_X1  g0804(.A1(new_n922), .A2(new_n706), .A3(new_n924), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT118), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n758), .A2(new_n310), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G87), .A2(new_n789), .B1(new_n752), .B2(G143), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n203), .B2(new_n754), .C1(new_n314), .C2(new_n756), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1007), .B(new_n1009), .C1(G50), .C2(new_n736), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n732), .A2(new_n253), .B1(new_n748), .B2(new_n340), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n722), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT116), .Z(new_n1015));
  OAI22_X1  g0815(.A1(new_n732), .A2(new_n737), .B1(new_n748), .B2(new_n755), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT52), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n735), .A2(new_n593), .B1(new_n744), .B2(new_n301), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n754), .A2(new_n741), .B1(new_n751), .B2(new_n966), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n275), .B1(new_n758), .B2(new_n245), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1017), .B(new_n1021), .C1(new_n971), .C2(new_n756), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT117), .Z(new_n1024));
  AOI21_X1  g0824(.A(new_n708), .B1(new_n1024), .B2(new_n728), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n729), .B1(new_n218), .B2(new_n213), .C1(new_n246), .C2(new_n952), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n954), .C2(new_n891), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1005), .A2(new_n1006), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1006), .B1(new_n1005), .B2(new_n1027), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n922), .A2(new_n924), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n915), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n925), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1031), .B1(new_n1034), .B2(new_n667), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G390));
  AOI22_X1  g0836(.A1(new_n736), .A2(G137), .B1(new_n733), .B2(G128), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n275), .B1(new_n759), .B2(G159), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n201), .C2(new_n744), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n754), .A2(new_n253), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT53), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT54), .B(G143), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n762), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n752), .A2(G125), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1039), .B(new_n1045), .C1(G132), .C2(new_n749), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G68), .A2(new_n789), .B1(new_n752), .B2(G294), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n218), .B2(new_n756), .C1(new_n245), .C2(new_n748), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n736), .A2(G107), .B1(new_n733), .B2(G283), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n553), .B2(new_n754), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1048), .A2(new_n1050), .A3(new_n269), .A4(new_n1007), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n728), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n806), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n248), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n708), .B(new_n1054), .C1(new_n871), .C2(new_n714), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n868), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n815), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n872), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n870), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n777), .A2(new_n322), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n701), .A2(new_n661), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1058), .B1(new_n1063), .B2(new_n867), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n861), .A2(new_n872), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(G330), .B(new_n778), .C1(new_n687), .C2(new_n692), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(new_n1058), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1061), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n871), .B2(new_n1059), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n844), .A2(G330), .A3(new_n778), .A4(new_n815), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1055), .B1(new_n1074), .B2(new_n706), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n864), .A2(new_n655), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n875), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1063), .A2(new_n867), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1069), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n844), .A2(G330), .A3(new_n778), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n815), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1068), .A2(new_n1058), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1072), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1083), .A2(KEYINPUT119), .A3(new_n868), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT119), .B1(new_n1083), .B2(new_n868), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1074), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n667), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1074), .B1(new_n1077), .B2(new_n1086), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1075), .B1(new_n1088), .B2(new_n1089), .ZN(G378));
  AND3_X1   g0890(.A1(new_n846), .A2(KEYINPUT102), .A3(new_n847), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT102), .B1(new_n846), .B2(new_n847), .ZN(new_n1092));
  OAI211_X1 g0892(.A(G330), .B(new_n862), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n299), .B1(new_n636), .B2(new_n637), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n268), .A3(new_n820), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n268), .A2(new_n820), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n299), .B(new_n1097), .C1(new_n636), .C2(new_n637), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT56), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT55), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT56), .B1(new_n1105), .B2(new_n1099), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1093), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n852), .A2(G330), .A3(new_n862), .A4(new_n1107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n873), .A2(KEYINPUT120), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1087), .A2(new_n1077), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT57), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT57), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1087), .B2(new_n1077), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1109), .A2(new_n1110), .A3(new_n873), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n873), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n667), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1107), .A2(new_n714), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n806), .A2(new_n201), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n748), .A2(new_n1126), .B1(new_n756), .B2(new_n947), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n761), .B2(new_n1042), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n736), .A2(G132), .B1(new_n733), .B2(G125), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n253), .C2(new_n758), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT59), .Z(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n752), .B2(G124), .ZN(new_n1132));
  AOI21_X1  g0932(.A(G33), .B1(new_n789), .B2(new_n765), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n744), .A2(new_n202), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n749), .A2(G107), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n752), .A2(G283), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n982), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n561), .B2(new_n762), .ZN(new_n1140));
  INV_X1    g0940(.A(G41), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n732), .A2(new_n245), .B1(new_n758), .B2(new_n203), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n722), .B(new_n1142), .C1(G97), .C2(new_n736), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT58), .ZN(new_n1145));
  AOI21_X1  g0945(.A(G41), .B1(new_n722), .B2(G33), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1134), .B(new_n1145), .C1(G50), .C2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n708), .B1(new_n1147), .B2(new_n728), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1124), .A2(new_n1125), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1114), .B2(new_n706), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1123), .A2(new_n1151), .ZN(G375));
  OR2_X1    g0952(.A1(new_n1086), .A2(new_n1077), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1086), .A2(new_n1077), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n907), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1086), .A2(new_n706), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT122), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n756), .A2(new_n253), .B1(new_n751), .B2(new_n1126), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1135), .B(new_n1159), .C1(G137), .C2(new_n749), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n733), .A2(G132), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n736), .A2(new_n1042), .B1(new_n759), .B2(G50), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n801), .B1(G159), .B2(new_n761), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n748), .A2(new_n741), .B1(new_n756), .B2(new_n301), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G97), .B2(new_n761), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n269), .B1(new_n736), .B2(G116), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n733), .A2(G294), .B1(new_n789), .B2(G77), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n987), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n751), .A2(new_n593), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1164), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1171), .A2(new_n728), .B1(new_n203), .B2(new_n806), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n707), .B(new_n1172), .C1(new_n815), .C2(new_n715), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1158), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1156), .A2(new_n1174), .ZN(G381));
  NOR4_X1   g0975(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1176));
  INV_X1    g0976(.A(G375), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(G381), .A2(G384), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT123), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n1075), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1182), .ZN(G407));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n650), .A3(new_n1182), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(G407), .A2(G213), .A3(new_n1184), .ZN(G409));
  NAND2_X1  g0985(.A1(new_n650), .A2(G213), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT125), .B1(new_n1086), .B2(new_n1077), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n668), .B1(new_n1187), .B2(KEYINPUT60), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n1154), .C1(KEYINPUT60), .C2(new_n1187), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1174), .A2(new_n1189), .A3(G384), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G384), .B1(new_n1174), .B2(new_n1189), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(G378), .B(new_n1151), .C1(new_n1116), .C2(new_n1122), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1111), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n907), .A3(new_n1198), .A4(new_n1115), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n706), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n1149), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT124), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1182), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1194), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1201), .B2(new_n1182), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1186), .B(new_n1193), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT62), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1186), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n650), .A2(G213), .A3(G2897), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1174), .A2(new_n1189), .ZN(new_n1212));
  INV_X1    g1012(.A(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1190), .A3(new_n1209), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1208), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT61), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1201), .A2(new_n1182), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT124), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1203), .A3(new_n1194), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT62), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1186), .A4(new_n1193), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1207), .A2(new_n1217), .A3(new_n1218), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n927), .A2(new_n955), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n1035), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(G393), .B(new_n773), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n959), .B2(G390), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT127), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1225), .B2(new_n1035), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(G390), .A2(KEYINPUT127), .A3(new_n955), .A4(new_n927), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1225), .A2(new_n1035), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1227), .B(KEYINPUT126), .Z(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1229), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1224), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT61), .B1(new_n1229), .B2(new_n1236), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1221), .A2(KEYINPUT63), .A3(new_n1186), .A4(new_n1193), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT63), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1208), .B2(new_n1216), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1206), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1239), .B(new_n1240), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1238), .A2(new_n1244), .ZN(G405));
  INV_X1    g1045(.A(new_n1193), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1182), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1194), .B(new_n1246), .C1(new_n1177), .C2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1123), .B2(new_n1151), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1194), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1193), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(new_n1237), .ZN(G402));
endmodule


