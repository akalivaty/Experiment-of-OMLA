

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(G543), .A2(G651), .ZN(n626) );
  XNOR2_X2 U550 ( .A(n516), .B(KEYINPUT65), .ZN(n735) );
  INV_X1 U551 ( .A(KEYINPUT27), .ZN(n610) );
  XNOR2_X1 U552 ( .A(n611), .B(n610), .ZN(n613) );
  NOR2_X1 U553 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U554 ( .A1(n679), .A2(n678), .ZN(n689) );
  NOR2_X1 U555 ( .A1(n691), .A2(n690), .ZN(n692) );
  INV_X1 U556 ( .A(KEYINPUT106), .ZN(n705) );
  INV_X1 U557 ( .A(G651), .ZN(n535) );
  NOR2_X1 U558 ( .A1(n538), .A2(G651), .ZN(n799) );
  NOR2_X1 U559 ( .A1(G2104), .A2(n517), .ZN(n878) );
  NOR2_X1 U560 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U561 ( .A(n760), .B(KEYINPUT109), .ZN(n761) );
  XNOR2_X1 U562 ( .A(n524), .B(KEYINPUT94), .ZN(G164) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X1 U564 ( .A(KEYINPUT66), .B(n514), .Z(n515) );
  XNOR2_X1 U565 ( .A(KEYINPUT17), .B(n515), .ZN(n592) );
  AND2_X1 U566 ( .A1(G138), .A2(n592), .ZN(n523) );
  INV_X1 U567 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n517), .A2(G2104), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n735), .A2(G102), .ZN(n521) );
  NAND2_X1 U570 ( .A1(G126), .A2(n878), .ZN(n519) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U572 ( .A1(G114), .A2(n879), .ZN(n518) );
  AND2_X1 U573 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n879), .A2(G113), .ZN(n526) );
  NAND2_X1 U577 ( .A1(G137), .A2(n592), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U579 ( .A1(G101), .A2(n735), .ZN(n527) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n527), .Z(n529) );
  NAND2_X1 U581 ( .A1(n878), .A2(G125), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n531), .A2(n530), .ZN(G160) );
  NAND2_X1 U584 ( .A1(G85), .A2(n626), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n538) );
  NOR2_X1 U586 ( .A1(n538), .A2(n535), .ZN(n794) );
  NAND2_X1 U587 ( .A1(G72), .A2(n794), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(KEYINPUT67), .B(n534), .ZN(n542) );
  NOR2_X1 U590 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n536), .Z(n537) );
  XNOR2_X2 U592 ( .A(KEYINPUT68), .B(n537), .ZN(n797) );
  NAND2_X1 U593 ( .A1(n797), .A2(G60), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n799), .A2(G47), .ZN(n539) );
  AND2_X1 U595 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(G290) );
  NAND2_X1 U597 ( .A1(G73), .A2(n794), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT2), .ZN(n550) );
  NAND2_X1 U599 ( .A1(n799), .A2(G48), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G61), .A2(n797), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n626), .A2(G86), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT86), .B(n546), .Z(n547) );
  NOR2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(G305) );
  XNOR2_X1 U606 ( .A(KEYINPUT80), .B(KEYINPUT7), .ZN(n562) );
  NAND2_X1 U607 ( .A1(n626), .A2(G89), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G76), .A2(n794), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n554), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G63), .A2(n797), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT79), .B(n555), .Z(n557) );
  NAND2_X1 U614 ( .A1(n799), .A2(G51), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U618 ( .A(n562), .B(n561), .ZN(G168) );
  XOR2_X1 U619 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U620 ( .A1(n799), .A2(G53), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G65), .A2(n797), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G91), .A2(n626), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G78), .A2(n794), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  OR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(G299) );
  NAND2_X1 U627 ( .A1(n799), .A2(G52), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G64), .A2(n797), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n626), .A2(G90), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT69), .B(n571), .Z(n573) );
  NAND2_X1 U632 ( .A1(n794), .A2(G77), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  NOR2_X1 U635 ( .A1(n576), .A2(n575), .ZN(G171) );
  NAND2_X1 U636 ( .A1(G50), .A2(n799), .ZN(n583) );
  NAND2_X1 U637 ( .A1(G75), .A2(n794), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G62), .A2(n797), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G88), .A2(n626), .ZN(n579) );
  XNOR2_X1 U641 ( .A(KEYINPUT87), .B(n579), .ZN(n580) );
  NOR2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U644 ( .A(n584), .B(KEYINPUT88), .ZN(G303) );
  NAND2_X1 U645 ( .A1(G49), .A2(n799), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G87), .A2(n538), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U648 ( .A1(n797), .A2(n587), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G74), .A2(G651), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT85), .B(n588), .Z(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(G288) );
  NOR2_X1 U652 ( .A1(G1384), .A2(G164), .ZN(n618) );
  AND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n615) );
  INV_X1 U654 ( .A(n615), .ZN(n591) );
  NOR2_X1 U655 ( .A1(n618), .A2(n591), .ZN(n756) );
  XOR2_X1 U656 ( .A(G2067), .B(KEYINPUT37), .Z(n753) );
  NAND2_X1 U657 ( .A1(n735), .A2(G104), .ZN(n595) );
  INV_X1 U658 ( .A(n592), .ZN(n593) );
  INV_X1 U659 ( .A(n593), .ZN(n882) );
  NAND2_X1 U660 ( .A1(G140), .A2(n882), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U662 ( .A(KEYINPUT34), .B(n596), .ZN(n603) );
  NAND2_X1 U663 ( .A1(n879), .A2(G116), .ZN(n597) );
  XNOR2_X1 U664 ( .A(KEYINPUT97), .B(n597), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n878), .A2(G128), .ZN(n598) );
  XOR2_X1 U666 ( .A(KEYINPUT96), .B(n598), .Z(n599) );
  NOR2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT35), .ZN(n602) );
  NOR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U670 ( .A(KEYINPUT36), .B(n604), .Z(n891) );
  AND2_X1 U671 ( .A1(n753), .A2(n891), .ZN(n927) );
  NAND2_X1 U672 ( .A1(n756), .A2(n927), .ZN(n752) );
  XNOR2_X1 U673 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U674 ( .A1(n968), .A2(n756), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT95), .B(n605), .Z(n606) );
  NAND2_X1 U676 ( .A1(n752), .A2(n606), .ZN(n725) );
  NAND2_X1 U677 ( .A1(n618), .A2(n615), .ZN(n680) );
  NAND2_X1 U678 ( .A1(G8), .A2(n680), .ZN(n718) );
  NOR2_X1 U679 ( .A1(G1981), .A2(G305), .ZN(n607) );
  XOR2_X1 U680 ( .A(n607), .B(KEYINPUT24), .Z(n608) );
  NOR2_X1 U681 ( .A1(n718), .A2(n608), .ZN(n723) );
  INV_X1 U682 ( .A(KEYINPUT100), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n680), .B(n609), .ZN(n638) );
  NAND2_X1 U684 ( .A1(G2072), .A2(n638), .ZN(n611) );
  INV_X1 U685 ( .A(n638), .ZN(n663) );
  NAND2_X1 U686 ( .A1(n663), .A2(G1956), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n656) );
  NAND2_X1 U688 ( .A1(G299), .A2(n656), .ZN(n614) );
  XOR2_X1 U689 ( .A(KEYINPUT28), .B(n614), .Z(n661) );
  XOR2_X1 U690 ( .A(G1996), .B(KEYINPUT102), .Z(n945) );
  INV_X1 U691 ( .A(n945), .ZN(n616) );
  AND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  AND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U694 ( .A(KEYINPUT26), .B(KEYINPUT103), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n680), .A2(G1341), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n636) );
  NAND2_X1 U698 ( .A1(G56), .A2(n797), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT14), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G43), .A2(n799), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n634) );
  NAND2_X1 U702 ( .A1(G81), .A2(n626), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT12), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT72), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n794), .A2(G68), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U707 ( .A(KEYINPUT13), .B(n631), .ZN(n632) );
  XNOR2_X1 U708 ( .A(KEYINPUT73), .B(n632), .ZN(n633) );
  XOR2_X2 U709 ( .A(KEYINPUT74), .B(n635), .Z(n981) );
  NOR2_X1 U710 ( .A1(n636), .A2(n981), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(KEYINPUT64), .ZN(n652) );
  NAND2_X1 U712 ( .A1(n638), .A2(G2067), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G1348), .A2(n680), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n653) );
  NAND2_X1 U715 ( .A1(G79), .A2(n794), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G54), .A2(n799), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(KEYINPUT76), .B(n643), .ZN(n647) );
  NAND2_X1 U719 ( .A1(G92), .A2(n626), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G66), .A2(n797), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U723 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT77), .B(n650), .Z(n895) );
  NOR2_X1 U726 ( .A1(n653), .A2(n895), .ZN(n651) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n655) );
  AND2_X1 U728 ( .A1(n895), .A2(n653), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n658) );
  NOR2_X1 U730 ( .A1(G299), .A2(n656), .ZN(n657) );
  NOR2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT104), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n662), .B(KEYINPUT29), .ZN(n670) );
  INV_X1 U734 ( .A(n663), .ZN(n664) );
  XNOR2_X1 U735 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U736 ( .A1(n664), .A2(n946), .ZN(n667) );
  INV_X1 U737 ( .A(G1961), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n665), .A2(n680), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n674) );
  AND2_X1 U740 ( .A1(n674), .A2(G171), .ZN(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT101), .B(n668), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n679) );
  NOR2_X1 U743 ( .A1(G1966), .A2(n718), .ZN(n691) );
  NOR2_X1 U744 ( .A1(G2084), .A2(n680), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n691), .A2(n688), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G8), .A2(n671), .ZN(n672) );
  XNOR2_X1 U747 ( .A(KEYINPUT30), .B(n672), .ZN(n673) );
  NOR2_X1 U748 ( .A1(G168), .A2(n673), .ZN(n676) );
  NOR2_X1 U749 ( .A1(G171), .A2(n674), .ZN(n675) );
  NOR2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT31), .B(n677), .Z(n678) );
  NAND2_X1 U752 ( .A1(G286), .A2(n689), .ZN(n685) );
  NOR2_X1 U753 ( .A1(G1971), .A2(n718), .ZN(n682) );
  NOR2_X1 U754 ( .A1(G2090), .A2(n680), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n683), .A2(G303), .ZN(n684) );
  NAND2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U758 ( .A1(n686), .A2(G8), .ZN(n687) );
  XNOR2_X1 U759 ( .A(n687), .B(KEYINPUT32), .ZN(n713) );
  NAND2_X1 U760 ( .A1(G8), .A2(n688), .ZN(n693) );
  INV_X1 U761 ( .A(n689), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n714) );
  INV_X1 U763 ( .A(KEYINPUT33), .ZN(n699) );
  NAND2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U765 ( .A(n718), .ZN(n694) );
  NAND2_X1 U766 ( .A1(n973), .A2(n694), .ZN(n695) );
  NAND2_X1 U767 ( .A1(n699), .A2(n695), .ZN(n697) );
  AND2_X1 U768 ( .A1(n714), .A2(n697), .ZN(n696) );
  NAND2_X1 U769 ( .A1(n713), .A2(n696), .ZN(n704) );
  INV_X1 U770 ( .A(n697), .ZN(n702) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n707) );
  NOR2_X1 U772 ( .A1(G303), .A2(G1971), .ZN(n698) );
  NOR2_X1 U773 ( .A1(n707), .A2(n698), .ZN(n970) );
  XOR2_X1 U774 ( .A(n970), .B(KEYINPUT105), .Z(n700) );
  AND2_X1 U775 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U776 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U778 ( .A(n706), .B(n705), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n707), .A2(KEYINPUT33), .ZN(n708) );
  NOR2_X1 U780 ( .A1(n718), .A2(n708), .ZN(n710) );
  XOR2_X1 U781 ( .A(G1981), .B(G305), .Z(n964) );
  INV_X1 U782 ( .A(n964), .ZN(n709) );
  NOR2_X1 U783 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n721) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n717) );
  NOR2_X1 U786 ( .A1(G2090), .A2(G303), .ZN(n715) );
  NAND2_X1 U787 ( .A1(G8), .A2(n715), .ZN(n716) );
  NAND2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n735), .A2(G95), .ZN(n727) );
  NAND2_X1 U794 ( .A1(G131), .A2(n882), .ZN(n726) );
  NAND2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U796 ( .A(KEYINPUT98), .B(n728), .Z(n732) );
  NAND2_X1 U797 ( .A1(G119), .A2(n878), .ZN(n730) );
  NAND2_X1 U798 ( .A1(G107), .A2(n879), .ZN(n729) );
  AND2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n888) );
  NAND2_X1 U801 ( .A1(G1991), .A2(n888), .ZN(n742) );
  NAND2_X1 U802 ( .A1(n878), .A2(G129), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G141), .A2(n882), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n738) );
  NAND2_X1 U805 ( .A1(n735), .A2(G105), .ZN(n736) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n736), .Z(n737) );
  NOR2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U808 ( .A1(n879), .A2(G117), .ZN(n739) );
  NAND2_X1 U809 ( .A1(n740), .A2(n739), .ZN(n875) );
  NAND2_X1 U810 ( .A1(G1996), .A2(n875), .ZN(n741) );
  NAND2_X1 U811 ( .A1(n742), .A2(n741), .ZN(n920) );
  AND2_X1 U812 ( .A1(n756), .A2(n920), .ZN(n748) );
  XNOR2_X1 U813 ( .A(KEYINPUT99), .B(n748), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n759) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n875), .ZN(n917) );
  NOR2_X1 U816 ( .A1(G1991), .A2(n888), .ZN(n923) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n745) );
  XOR2_X1 U818 ( .A(n745), .B(KEYINPUT107), .Z(n746) );
  NOR2_X1 U819 ( .A1(n923), .A2(n746), .ZN(n747) );
  NOR2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U821 ( .A1(n917), .A2(n749), .ZN(n750) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n750), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n755) );
  NOR2_X1 U824 ( .A1(n753), .A2(n891), .ZN(n754) );
  XOR2_X1 U825 ( .A(KEYINPUT108), .B(n754), .Z(n935) );
  NAND2_X1 U826 ( .A1(n755), .A2(n935), .ZN(n757) );
  NAND2_X1 U827 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U828 ( .A1(n759), .A2(n758), .ZN(n762) );
  XOR2_X1 U829 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n760) );
  XNOR2_X1 U830 ( .A(n762), .B(n761), .ZN(G329) );
  INV_X1 U831 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U832 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U833 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  NAND2_X1 U835 ( .A1(G108), .A2(G120), .ZN(n763) );
  NOR2_X1 U836 ( .A1(G237), .A2(n763), .ZN(n764) );
  NAND2_X1 U837 ( .A1(G69), .A2(n764), .ZN(n833) );
  NAND2_X1 U838 ( .A1(n833), .A2(G567), .ZN(n769) );
  NOR2_X1 U839 ( .A1(G220), .A2(G219), .ZN(n765) );
  XOR2_X1 U840 ( .A(KEYINPUT22), .B(n765), .Z(n766) );
  NOR2_X1 U841 ( .A1(G218), .A2(n766), .ZN(n767) );
  NAND2_X1 U842 ( .A1(G96), .A2(n767), .ZN(n834) );
  NAND2_X1 U843 ( .A1(n834), .A2(G2106), .ZN(n768) );
  AND2_X1 U844 ( .A1(n769), .A2(n768), .ZN(G319) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  XNOR2_X1 U846 ( .A(G860), .B(KEYINPUT75), .ZN(n778) );
  OR2_X1 U847 ( .A1(n981), .A2(n778), .ZN(G153) );
  XOR2_X1 U848 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n771) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U850 ( .A(n771), .B(n770), .ZN(G223) );
  INV_X1 U851 ( .A(G223), .ZN(n828) );
  NAND2_X1 U852 ( .A1(n828), .A2(G567), .ZN(n772) );
  XOR2_X1 U853 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U854 ( .A(G171), .ZN(G301) );
  NOR2_X1 U855 ( .A1(n895), .A2(G868), .ZN(n774) );
  INV_X1 U856 ( .A(G868), .ZN(n806) );
  NOR2_X1 U857 ( .A1(n806), .A2(G301), .ZN(n773) );
  NOR2_X1 U858 ( .A1(n774), .A2(n773), .ZN(G284) );
  NAND2_X1 U859 ( .A1(G299), .A2(n806), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G868), .A2(G286), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U862 ( .A(KEYINPUT81), .B(n777), .Z(G297) );
  NAND2_X1 U863 ( .A1(n778), .A2(G559), .ZN(n779) );
  INV_X1 U864 ( .A(n895), .ZN(n975) );
  NAND2_X1 U865 ( .A1(n779), .A2(n975), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT82), .ZN(n781) );
  XNOR2_X1 U867 ( .A(KEYINPUT16), .B(n781), .ZN(G148) );
  NOR2_X1 U868 ( .A1(n981), .A2(G868), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n975), .A2(G868), .ZN(n782) );
  NOR2_X1 U870 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U872 ( .A1(G99), .A2(n735), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G111), .A2(n879), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n878), .A2(G123), .ZN(n787) );
  XOR2_X1 U876 ( .A(KEYINPUT18), .B(n787), .Z(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G135), .A2(n882), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n924) );
  XOR2_X1 U880 ( .A(n924), .B(G2096), .Z(n793) );
  XNOR2_X1 U881 ( .A(G2100), .B(KEYINPUT83), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(G156) );
  NAND2_X1 U883 ( .A1(G93), .A2(n626), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G80), .A2(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n803) );
  NAND2_X1 U886 ( .A1(G67), .A2(n797), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT84), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G559), .A2(n975), .ZN(n815) );
  XNOR2_X1 U892 ( .A(n981), .B(n815), .ZN(n804) );
  NOR2_X1 U893 ( .A1(G860), .A2(n804), .ZN(n805) );
  XOR2_X1 U894 ( .A(n807), .B(n805), .Z(G145) );
  INV_X1 U895 ( .A(G303), .ZN(G166) );
  NAND2_X1 U896 ( .A1(n806), .A2(n807), .ZN(n818) );
  XNOR2_X1 U897 ( .A(G299), .B(G305), .ZN(n814) );
  XNOR2_X1 U898 ( .A(KEYINPUT89), .B(KEYINPUT19), .ZN(n808) );
  XOR2_X1 U899 ( .A(n808), .B(n807), .Z(n811) );
  XNOR2_X1 U900 ( .A(n981), .B(G290), .ZN(n809) );
  XNOR2_X1 U901 ( .A(n809), .B(G166), .ZN(n810) );
  XNOR2_X1 U902 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n812), .B(G288), .ZN(n813) );
  XNOR2_X1 U904 ( .A(n814), .B(n813), .ZN(n896) );
  XNOR2_X1 U905 ( .A(n896), .B(n815), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n816), .A2(G868), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U908 ( .A(n819), .B(KEYINPUT90), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2078), .A2(G2084), .ZN(n820) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U911 ( .A1(G2090), .A2(n821), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n822) );
  XNOR2_X1 U913 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G2072), .A2(n824), .ZN(G158) );
  NAND2_X1 U915 ( .A1(G661), .A2(G483), .ZN(n825) );
  XOR2_X1 U916 ( .A(KEYINPUT92), .B(n825), .Z(n826) );
  NAND2_X1 U917 ( .A1(n826), .A2(G319), .ZN(n827) );
  XNOR2_X1 U918 ( .A(n827), .B(KEYINPUT93), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U922 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT111), .B(n832), .Z(G188) );
  XOR2_X1 U926 ( .A(G120), .B(KEYINPUT112), .Z(G236) );
  NOR2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G325) );
  XNOR2_X1 U928 ( .A(KEYINPUT113), .B(G325), .ZN(G261) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  XOR2_X1 U932 ( .A(G1981), .B(G1966), .Z(n836) );
  XNOR2_X1 U933 ( .A(G1991), .B(G1996), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n846) );
  XOR2_X1 U935 ( .A(KEYINPUT115), .B(KEYINPUT117), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1956), .B(G2474), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1961), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT41), .B(KEYINPUT116), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(G229) );
  XOR2_X1 U945 ( .A(G2100), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2072), .B(KEYINPUT42), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n849), .B(G2678), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2090), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(KEYINPUT114), .B(G2096), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U955 ( .A1(n878), .A2(G124), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G112), .A2(n879), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n735), .A2(G100), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G136), .A2(n882), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(G162) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n864) );
  XNOR2_X1 U964 ( .A(G164), .B(KEYINPUT118), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n874) );
  NAND2_X1 U966 ( .A1(n735), .A2(G103), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G139), .A2(n882), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G127), .A2(n878), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G115), .A2(n879), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n931) );
  XOR2_X1 U974 ( .A(n931), .B(G162), .Z(n872) );
  XNOR2_X1 U975 ( .A(n924), .B(n872), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n875), .B(G160), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n893) );
  NAND2_X1 U979 ( .A1(G130), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n887) );
  NAND2_X1 U982 ( .A1(n735), .A2(G106), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n891), .B(n890), .Z(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U990 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n895), .B(G286), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n898), .B(G171), .ZN(n899) );
  NOR2_X1 U994 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2451), .B(G2430), .Z(n901) );
  XNOR2_X1 U996 ( .A(G2438), .B(G2443), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n907) );
  XOR2_X1 U998 ( .A(G2435), .B(G2454), .Z(n903) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1001 ( .A(G2446), .B(G2427), .Z(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n907), .B(n906), .Z(n908) );
  NAND2_X1 U1004 ( .A1(G14), .A2(n908), .ZN(n914) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  INV_X1 U1013 ( .A(n914), .ZN(G401) );
  XNOR2_X1 U1014 ( .A(G2090), .B(G162), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n915), .B(KEYINPUT121), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT51), .B(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n930) );
  XNOR2_X1 U1019 ( .A(G160), .B(G2084), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n921), .B(KEYINPUT119), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n928), .B(KEYINPUT120), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n938) );
  XOR2_X1 U1026 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n934), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n960) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n960), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n955) );
  XOR2_X1 U1037 ( .A(G1991), .B(G25), .Z(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(G2067), .B(G26), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n950) );
  XOR2_X1 U1042 ( .A(n945), .B(G32), .Z(n948) );
  XOR2_X1 U1043 ( .A(n946), .B(G27), .Z(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1049 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n960), .B(n959), .ZN(n962) );
  INV_X1 U1053 ( .A(G29), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n963), .ZN(n1018) );
  XNOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .ZN(n988) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT57), .B(n966), .ZN(n986) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G301), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n980) );
  NAND2_X1 U1062 ( .A1(G303), .A2(G1971), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G299), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n978) );
  XOR2_X1 U1067 ( .A(G1348), .B(n975), .Z(n976) );
  XNOR2_X1 U1068 ( .A(KEYINPUT122), .B(n976), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n981), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1073 ( .A(KEYINPUT123), .B(n984), .Z(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n1016) );
  INV_X1 U1076 ( .A(G16), .ZN(n1014) );
  XOR2_X1 U1077 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n995) );
  XNOR2_X1 U1078 ( .A(G1986), .B(G24), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1081 ( .A(G1976), .B(KEYINPUT126), .Z(n991) );
  XNOR2_X1 U1082 ( .A(G23), .B(n991), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n1011) );
  XOR2_X1 U1085 ( .A(G1966), .B(G21), .Z(n1006) );
  XOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .Z(n996) );
  XNOR2_X1 U1087 ( .A(G4), .B(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G6), .B(G1981), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G20), .B(G1956), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT124), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(KEYINPUT60), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G5), .B(G1961), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT125), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

