//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n214), .B1(new_n202), .B2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n217), .A2(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n216), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT65), .B(G238), .Z(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n213), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n211), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G13), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n213), .A2(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n223), .B(new_n235), .C1(new_n220), .C2(new_n225), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT0), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n233), .B(new_n237), .C1(new_n232), .C2(new_n231), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(G223), .B1(new_n265), .B2(G77), .ZN(new_n266));
  INV_X1    g0066(.A(G222), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n261), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n257), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n208), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G33), .A3(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(new_n271), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n208), .B1(KEYINPUT68), .B2(new_n272), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT69), .A3(new_n279), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n276), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n282), .B2(new_n284), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n275), .B(new_n289), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT74), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n299), .A2(KEYINPUT70), .A3(new_n208), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT70), .B1(new_n299), .B2(new_n208), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n234), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OR3_X1    g0105(.A1(new_n302), .A2(KEYINPUT71), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT71), .B1(new_n302), .B2(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(G50), .C1(G1), .C2(new_n209), .ZN(new_n309));
  OAI21_X1  g0109(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n310));
  INV_X1    g0110(.A(G150), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G20), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n259), .A2(G20), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n310), .B1(new_n311), .B2(new_n313), .C1(new_n314), .C2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n302), .B1(new_n201), .B2(new_n305), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT9), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT9), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n320), .A2(KEYINPUT73), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT73), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n295), .B(new_n298), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n297), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n295), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT10), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n293), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n319), .B(new_n330), .C1(G179), .C2(new_n293), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n312), .A2(G50), .B1(G20), .B2(new_n229), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n316), .B2(new_n217), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n302), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT11), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n305), .A2(new_n229), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n209), .A2(G1), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n302), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G68), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n336), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n291), .A2(G238), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT75), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n269), .B2(new_n290), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G232), .B2(new_n262), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n289), .B(new_n343), .C1(new_n347), .C2(new_n273), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT13), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n349), .B2(new_n296), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g0156(.A(new_n342), .B(KEYINPUT76), .Z(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT14), .B1(new_n353), .B2(new_n329), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n349), .A2(new_n359), .A3(G169), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(G179), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n356), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n291), .A2(G232), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n289), .A2(new_n366), .A3(new_n296), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT80), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n369), .B(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(G223), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n372));
  OAI211_X1 g0172(.A(G226), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n274), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT81), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n377), .A3(new_n274), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n289), .A2(new_n366), .A3(new_n375), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n368), .A2(new_n380), .B1(new_n381), .B2(new_n354), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n314), .A2(new_n339), .ZN(new_n383));
  XOR2_X1   g0183(.A(new_n383), .B(KEYINPUT79), .Z(new_n384));
  AOI22_X1  g0184(.A1(new_n308), .A2(new_n384), .B1(new_n305), .B2(new_n314), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n202), .A2(new_n229), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G58), .A2(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n312), .A2(G159), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n268), .A2(new_n392), .A3(G20), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT77), .B1(new_n263), .B2(new_n264), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n260), .A2(new_n395), .A3(new_n261), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n396), .A3(new_n209), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n391), .C1(new_n398), .C2(new_n229), .ZN(new_n399));
  XOR2_X1   g0199(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n400));
  OAI21_X1  g0200(.A(new_n392), .B1(new_n268), .B2(G20), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n229), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n403), .B2(new_n390), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n302), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n385), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n365), .B1(new_n382), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n289), .A2(new_n366), .A3(new_n375), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n408), .A2(G200), .B1(new_n367), .B2(new_n379), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n385), .A4(new_n405), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G179), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n289), .A2(new_n366), .A3(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n380), .B1(new_n381), .B2(new_n329), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n414), .A2(new_n406), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n414), .B2(new_n406), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT82), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n406), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT82), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n414), .A2(new_n406), .A3(new_n415), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n411), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n426), .A2(new_n316), .B1(new_n209), .B2(new_n217), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n314), .A2(new_n313), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n302), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n340), .A2(G77), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(G77), .C2(new_n304), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n265), .A2(G107), .ZN(new_n432));
  INV_X1    g0232(.A(new_n262), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n432), .B1(new_n269), .B2(new_n215), .C1(new_n228), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n274), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n289), .C1(new_n218), .C2(new_n292), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n436), .B2(G200), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n296), .B2(new_n436), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n329), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n431), .C1(G179), .C2(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT72), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n332), .A2(new_n364), .A3(new_n425), .A4(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n268), .A2(new_n209), .A3(G87), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT22), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n209), .B2(G107), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G116), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n447), .A2(new_n448), .B1(new_n450), .B2(new_n209), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT24), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n302), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n305), .A2(new_n224), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT25), .ZN(new_n456));
  OAI221_X1 g0256(.A(new_n304), .B1(G1), .B2(new_n259), .C1(new_n300), .C2(new_n301), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(G107), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n282), .A2(new_n284), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n286), .A2(G45), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(G274), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n465), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT69), .B1(new_n283), .B2(new_n279), .ZN(new_n468));
  AND4_X1   g0268(.A1(KEYINPUT69), .A2(new_n277), .A3(new_n279), .A4(new_n271), .ZN(new_n469));
  OAI211_X1 g0269(.A(G264), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT91), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n461), .A2(new_n472), .A3(G264), .A4(new_n467), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n262), .A2(G257), .B1(G33), .B2(G294), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n268), .A2(G250), .A3(new_n257), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n273), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT92), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT92), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n480), .B(new_n477), .C1(new_n471), .C2(new_n473), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n466), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n354), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n466), .A3(new_n470), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(KEYINPUT90), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(KEYINPUT90), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n296), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n460), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G179), .B(new_n466), .C1(new_n479), .C2(new_n481), .ZN(new_n490));
  OAI21_X1  g0290(.A(G169), .B1(new_n485), .B2(new_n486), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n491), .B1(new_n454), .B2(new_n459), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT93), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n460), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT93), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n482), .A2(new_n354), .B1(new_n487), .B2(new_n296), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n460), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n462), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n223), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n461), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(G274), .B(new_n499), .C1(new_n468), .C2(new_n469), .ZN(new_n502));
  OAI211_X1 g0302(.A(G238), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n449), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n274), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT19), .B1(new_n315), .B2(G97), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n268), .A2(new_n209), .A3(G68), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(KEYINPUT87), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n268), .A2(new_n513), .A3(new_n209), .A4(G68), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT75), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n344), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT19), .ZN(new_n518));
  NOR2_X1   g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n518), .A2(new_n209), .B1(new_n222), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n302), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n426), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n304), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n458), .A2(G87), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT88), .B1(new_n509), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n518), .A2(new_n209), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(new_n222), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n514), .A3(new_n512), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n523), .B1(new_n531), .B2(new_n302), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT88), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n508), .A4(new_n525), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G190), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n527), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n521), .B(new_n524), .C1(new_n426), .C2(new_n457), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n507), .A2(G169), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT86), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n461), .A2(new_n500), .B1(new_n505), .B2(new_n274), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G179), .A3(new_n502), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n539), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n305), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n457), .B2(G97), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  OR2_X1    g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT85), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n262), .A2(G250), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n554), .A2(new_n555), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n268), .A2(G244), .A3(new_n257), .A4(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n554), .A2(new_n555), .B1(G33), .B2(G283), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n556), .A2(new_n557), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n274), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n465), .B1(new_n282), .B2(new_n284), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G257), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n466), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G190), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n401), .A2(new_n402), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n219), .A2(new_n224), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n519), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n572), .B2(KEYINPUT6), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n312), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n568), .B1(new_n567), .B2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n302), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n562), .A2(new_n466), .A3(new_n564), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n552), .A2(new_n566), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n565), .A2(new_n412), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n329), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n550), .A2(new_n551), .ZN(new_n583));
  INV_X1    g0383(.A(new_n302), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n569), .A2(new_n574), .ZN(new_n585));
  INV_X1    g0385(.A(new_n576), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G283), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n590), .B(new_n209), .C1(G33), .C2(new_n219), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n299), .A2(new_n208), .ZN(new_n592));
  INV_X1    g0392(.A(G116), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g0395(.A(new_n595), .B(KEYINPUT20), .Z(new_n596));
  NAND3_X1  g0396(.A1(new_n303), .A2(G20), .A3(new_n593), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n593), .C2(new_n457), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n461), .A2(G270), .A3(new_n467), .ZN(new_n600));
  OAI211_X1 g0400(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n260), .A2(G303), .A3(new_n261), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n604), .A2(KEYINPUT89), .A3(new_n274), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT89), .B1(new_n604), .B2(new_n274), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n466), .B(new_n600), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G200), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n599), .B(new_n608), .C1(new_n296), .C2(new_n607), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n598), .A2(G169), .A3(new_n607), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n598), .A2(new_n607), .A3(KEYINPUT21), .A4(G169), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n607), .A2(new_n412), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n598), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n609), .A2(new_n612), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n546), .A2(new_n589), .A3(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n443), .A2(new_n493), .A3(new_n498), .A4(new_n617), .ZN(G372));
  NAND4_X1  g0418(.A1(new_n532), .A2(new_n536), .A3(new_n508), .A4(new_n525), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n539), .A2(new_n542), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n538), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n622), .A2(new_n588), .A3(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(new_n588), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n537), .A3(new_n545), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n625), .B2(KEYINPUT26), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n495), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n580), .A2(new_n588), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n619), .C1(new_n497), .C2(new_n460), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n626), .B(new_n621), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n443), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n356), .A2(new_n440), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n362), .A2(new_n357), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n411), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n416), .A2(new_n417), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n328), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n633), .A2(new_n331), .A3(new_n639), .ZN(G369));
  INV_X1    g0440(.A(new_n303), .ZN(new_n641));
  OR3_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .A3(G20), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT27), .B1(new_n641), .B2(G20), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n460), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n493), .A2(new_n498), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n492), .A2(new_n646), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n627), .ZN(new_n651));
  INV_X1    g0451(.A(new_n646), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n599), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n616), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n492), .A2(new_n652), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n627), .A2(new_n646), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n493), .A2(new_n498), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(G399));
  NOR2_X1   g0462(.A1(new_n235), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n529), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n664), .A2(new_n206), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(KEYINPUT94), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(KEYINPUT94), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n493), .A2(new_n498), .A3(new_n617), .A4(new_n652), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT31), .ZN(new_n673));
  AOI21_X1  g0473(.A(G179), .B1(new_n541), .B2(new_n502), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n607), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT95), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n607), .A3(KEYINPUT95), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n565), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n482), .ZN(new_n680));
  INV_X1    g0480(.A(new_n473), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n472), .B1(new_n563), .B2(G264), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n478), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n480), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n474), .A2(KEYINPUT92), .A3(new_n478), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n535), .A2(new_n466), .A3(new_n564), .A4(new_n562), .ZN(new_n687));
  INV_X1    g0487(.A(new_n606), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n604), .A2(KEYINPUT89), .A3(new_n274), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(G179), .A3(new_n466), .A4(new_n600), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT30), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n680), .B1(new_n693), .B2(KEYINPUT96), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT96), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n479), .A2(new_n481), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n614), .A2(new_n535), .A3(new_n565), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n686), .A2(new_n692), .A3(KEYINPUT30), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT97), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n697), .A2(new_n698), .A3(new_n696), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT96), .B1(new_n703), .B2(new_n693), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n699), .A2(new_n695), .B1(new_n482), .B2(new_n679), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT97), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n707), .A3(new_n646), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n673), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n703), .A2(new_n693), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n680), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n671), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n632), .A2(new_n715), .A3(new_n652), .ZN(new_n716));
  INV_X1    g0516(.A(new_n621), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n630), .A2(new_n619), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n489), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n719), .B2(new_n628), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n622), .A2(new_n588), .ZN(new_n721));
  MUX2_X1   g0521(.A(new_n625), .B(new_n721), .S(KEYINPUT26), .Z(new_n722));
  AOI21_X1  g0522(.A(new_n646), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n716), .B1(new_n723), .B2(new_n715), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n670), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR2_X1   g0526(.A1(new_n234), .A2(G20), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G45), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n664), .A2(G1), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n657), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n655), .ZN(new_n732));
  INV_X1    g0532(.A(new_n235), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G355), .A3(new_n268), .ZN(new_n734));
  INV_X1    g0534(.A(G45), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n251), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n394), .A2(new_n396), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n235), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G45), .B2(new_n206), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n734), .B1(G116), .B2(new_n733), .C1(new_n736), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n208), .B1(G20), .B2(new_n329), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT33), .B(G317), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n412), .A2(new_n354), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n209), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n412), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n749), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n747), .A2(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(new_n296), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n748), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n268), .B(new_n754), .C1(G326), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G294), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n209), .B1(new_n760), .B2(G190), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G303), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n354), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n755), .A2(new_n751), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n763), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n749), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n749), .A2(new_n760), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n762), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n750), .A2(new_n229), .B1(new_n752), .B2(new_n217), .ZN(new_n778));
  INV_X1    g0578(.A(new_n766), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n265), .B(new_n778), .C1(G58), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n761), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n771), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n756), .A2(new_n201), .B1(new_n769), .B2(new_n224), .ZN(new_n786));
  INV_X1    g0586(.A(new_n765), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(G87), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n780), .A2(new_n782), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n776), .A2(new_n777), .A3(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n729), .B(new_n746), .C1(new_n790), .C2(new_n744), .ZN(new_n791));
  INV_X1    g0591(.A(new_n743), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n655), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n732), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  INV_X1    g0595(.A(new_n714), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n431), .A2(new_n646), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n438), .A2(new_n440), .A3(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT99), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n440), .A2(new_n652), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n632), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n646), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n632), .A2(new_n652), .A3(new_n801), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n730), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n796), .B2(new_n807), .ZN(new_n809));
  INV_X1    g0609(.A(new_n744), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n756), .A2(new_n811), .B1(new_n750), .B2(new_n311), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n766), .A2(new_n813), .B1(new_n752), .B2(new_n783), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n769), .A2(new_n229), .B1(new_n771), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G50), .B2(new_n787), .ZN(new_n820));
  INV_X1    g0620(.A(new_n737), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G58), .B2(new_n781), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n816), .A2(new_n817), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n769), .A2(new_n222), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n750), .A2(new_n770), .B1(new_n752), .B2(new_n593), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(G107), .C2(new_n787), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n756), .A2(new_n763), .B1(new_n771), .B2(new_n753), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n268), .B(new_n827), .C1(G294), .C2(new_n779), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n828), .A3(new_n782), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n810), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n744), .A2(new_n741), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n729), .B(new_n830), .C1(new_n217), .C2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n799), .B(new_n800), .C1(new_n440), .C2(new_n652), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n742), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n809), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  NOR2_X1   g0636(.A1(new_n727), .A2(new_n286), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n357), .A2(new_n646), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n363), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n357), .B(new_n646), .C1(new_n362), .C2(new_n356), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n803), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT40), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n409), .A2(new_n385), .A3(new_n405), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n308), .A2(new_n384), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n305), .A2(new_n314), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n391), .B1(new_n398), .B2(new_n229), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT100), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT100), .B(new_n391), .C1(new_n398), .C2(new_n229), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n400), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n399), .A2(new_n302), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n843), .B1(new_n853), .B2(new_n644), .ZN(new_n854));
  INV_X1    g0654(.A(new_n414), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n644), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n406), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n843), .A2(new_n419), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n853), .A2(new_n644), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n862), .B(KEYINPUT38), .C1(new_n424), .C2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n843), .A2(new_n419), .A3(new_n859), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(new_n860), .ZN(new_n867));
  INV_X1    g0667(.A(new_n411), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n859), .B1(new_n868), .B2(new_n637), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n842), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n707), .A2(new_n646), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n702), .A2(new_n872), .B1(new_n672), .B2(KEYINPUT31), .ZN(new_n873));
  AND4_X1   g0673(.A1(KEYINPUT31), .A2(new_n702), .A3(new_n646), .A4(new_n707), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n841), .B(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT101), .ZN(new_n876));
  INV_X1    g0676(.A(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n709), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT101), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n841), .A4(new_n871), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n862), .B1(new_n424), .B2(new_n863), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n865), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n864), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n883), .A3(new_n841), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n876), .A2(new_n880), .B1(new_n842), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n878), .A2(new_n443), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n887), .A2(new_n888), .A3(new_n671), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n864), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n362), .A2(new_n357), .A3(new_n652), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT39), .B1(new_n864), .B2(new_n870), .ZN(new_n893));
  OR3_X1    g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n356), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n635), .A2(new_n895), .A3(new_n838), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n838), .B1(new_n635), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n440), .A2(new_n646), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n806), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n901), .A2(new_n883), .B1(new_n638), .B2(new_n644), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n639), .A2(new_n331), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n724), .B2(new_n443), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n903), .B(new_n905), .Z(new_n906));
  AOI21_X1  g0706(.A(new_n837), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n890), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(G116), .A3(new_n210), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n386), .A2(new_n206), .A3(new_n217), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n229), .A2(G50), .ZN(new_n914));
  OAI211_X1 g0714(.A(G1), .B(new_n234), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT102), .Z(G367));
  INV_X1    g0717(.A(new_n738), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n745), .B1(new_n733), .B2(new_n426), .C1(new_n918), .C2(new_n246), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n919), .A2(new_n730), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n821), .B1(new_n770), .B2(new_n752), .C1(new_n759), .C2(new_n750), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT46), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n765), .B2(new_n593), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n922), .B(new_n924), .C1(new_n224), .C2(new_n761), .ZN(new_n925));
  INV_X1    g0725(.A(new_n769), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(G97), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n763), .B2(new_n766), .ZN(new_n928));
  XNOR2_X1  g0728(.A(KEYINPUT108), .B(G311), .ZN(new_n929));
  INV_X1    g0729(.A(G317), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n756), .A2(new_n929), .B1(new_n771), .B2(new_n930), .ZN(new_n931));
  NOR4_X1   g0731(.A1(new_n921), .A2(new_n925), .A3(new_n928), .A4(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n771), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n757), .A2(G143), .B1(new_n933), .B2(G137), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(new_n201), .B2(new_n752), .C1(new_n783), .C2(new_n750), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n761), .A2(new_n229), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n202), .A2(new_n765), .B1(new_n766), .B2(new_n311), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n265), .B1(new_n926), .B2(G77), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT109), .Z(new_n940));
  AOI21_X1  g0740(.A(new_n932), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT47), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n652), .B1(new_n532), .B2(new_n525), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n717), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT103), .Z(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n622), .B2(new_n943), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n920), .B1(new_n810), .B2(new_n942), .C1(new_n946), .C2(new_n792), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT110), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n663), .B(KEYINPUT41), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n661), .A2(new_n659), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n646), .B1(new_n583), .B2(new_n587), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n630), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n624), .A2(new_n646), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT44), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n954), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n661), .A2(new_n958), .A3(new_n659), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n957), .A2(new_n658), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n961), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n657), .B(new_n650), .C1(new_n963), .C2(new_n956), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n650), .A2(KEYINPUT107), .A3(new_n660), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT107), .B1(new_n650), .B2(new_n660), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n661), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n657), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n656), .A3(new_n661), .A4(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n962), .A2(new_n964), .A3(new_n970), .A4(new_n725), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n949), .B1(new_n971), .B2(new_n725), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n728), .A2(G1), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n661), .A2(new_n954), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n630), .A2(new_n492), .A3(new_n951), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n646), .B1(new_n977), .B2(new_n588), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n975), .B2(KEYINPUT42), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n976), .A2(new_n979), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT104), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT104), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n980), .A2(new_n984), .A3(KEYINPUT105), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n658), .A2(new_n954), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT105), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n982), .A2(new_n987), .A3(new_n983), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n987), .B1(new_n982), .B2(new_n983), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n980), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n985), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n986), .B1(new_n985), .B2(new_n990), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n948), .B1(new_n974), .B2(new_n993), .ZN(G387));
  OR2_X1    g0794(.A1(new_n970), .A2(new_n725), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n664), .B1(new_n970), .B2(new_n725), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n648), .A2(new_n649), .A3(new_n743), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n756), .A2(new_n767), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n750), .A2(new_n929), .B1(new_n752), .B2(new_n763), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G317), .C2(new_n779), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT48), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(KEYINPUT48), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n787), .A2(G294), .B1(new_n781), .B2(G283), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G116), .A2(new_n926), .B1(new_n933), .B2(G326), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n821), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n750), .A2(new_n314), .B1(new_n752), .B2(new_n229), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n787), .A2(G77), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n771), .B2(new_n311), .C1(new_n783), .C2(new_n756), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n779), .A2(G50), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n781), .A2(new_n522), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1014), .A2(new_n927), .A3(new_n737), .A4(new_n1015), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1011), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n810), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n243), .A2(G45), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n918), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n235), .A2(new_n265), .A3(new_n665), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n314), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT50), .B1(new_n314), .B2(G50), .ZN(new_n1023));
  AOI21_X1  g0823(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n665), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1020), .A2(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n733), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n729), .B(new_n1018), .C1(new_n745), .C2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n995), .A2(new_n996), .B1(new_n997), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n973), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n968), .B2(new_n969), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT111), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(G393));
  NAND3_X1  g0833(.A1(new_n962), .A2(new_n964), .A3(new_n973), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n918), .A2(new_n255), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n745), .B1(new_n733), .B2(new_n219), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n730), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT113), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n824), .B(new_n821), .C1(G143), .C2(new_n933), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n756), .A2(new_n311), .B1(new_n766), .B2(new_n783), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n750), .A2(new_n201), .B1(new_n752), .B2(new_n314), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G68), .B2(new_n787), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n781), .A2(G77), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n265), .B1(new_n769), .B2(new_n224), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n765), .A2(new_n770), .B1(new_n771), .B2(new_n767), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n752), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1047), .C1(G294), .C2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n756), .A2(new_n930), .B1(new_n766), .B2(new_n753), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n750), .A2(new_n763), .B1(new_n761), .B2(new_n593), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT114), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1045), .A2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1038), .B1(new_n810), .B2(new_n1055), .C1(new_n958), .C2(new_n792), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n971), .A2(new_n663), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n964), .A2(new_n962), .B1(new_n970), .B2(new_n725), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1034), .B(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(KEYINPUT115), .ZN(new_n1060));
  OAI211_X1 g0860(.A(G330), .B(new_n833), .C1(new_n873), .C2(new_n712), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n833), .B1(new_n896), .B2(new_n897), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n709), .B2(new_n877), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1061), .A2(new_n898), .B1(new_n1063), .B2(G330), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n806), .A2(new_n900), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1060), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n898), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n714), .B2(new_n833), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n874), .B1(new_n673), .B2(new_n708), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1070), .A2(new_n671), .A3(new_n1062), .ZN(new_n1071));
  OAI211_X1 g0871(.A(KEYINPUT115), .B(new_n1065), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n899), .B1(new_n723), .B2(new_n801), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1061), .B2(new_n898), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n671), .B1(new_n709), .B2(new_n877), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1068), .B1(new_n1076), .B2(new_n833), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n864), .A2(new_n870), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n892), .B(new_n1081), .C1(new_n1074), .C2(new_n898), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n892), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n901), .A2(new_n1083), .B1(new_n891), .B2(new_n893), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n714), .A2(new_n833), .A3(new_n1068), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1071), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1076), .A2(new_n443), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n905), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1080), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1078), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1089), .B1(new_n1095), .B2(new_n1092), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n663), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n741), .B1(new_n891), .B2(new_n893), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n224), .A2(new_n750), .B1(new_n766), .B2(new_n593), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n752), .A2(new_n219), .B1(new_n771), .B2(new_n759), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n268), .B1(new_n787), .B2(G87), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G283), .A2(new_n757), .B1(new_n926), .B2(G68), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n1044), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n756), .A2(new_n1105), .B1(new_n750), .B2(new_n811), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G132), .B2(new_n779), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n268), .B1(new_n769), .B2(new_n201), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n765), .A2(new_n311), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT53), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1112), .A2(new_n1113), .B1(G159), .B2(new_n781), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n752), .A2(new_n1115), .B1(new_n771), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1114), .B(new_n1118), .C1(new_n1113), .C2(new_n1112), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1104), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n744), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n729), .B1(new_n314), .B2(new_n831), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1098), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1090), .B2(new_n973), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1097), .A2(new_n1124), .ZN(G378));
  INV_X1    g0925(.A(KEYINPUT118), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n884), .A2(new_n842), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n879), .B1(new_n1063), .B2(new_n871), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1081), .A2(KEYINPUT40), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1070), .A2(new_n1129), .A3(KEYINPUT101), .A4(new_n1062), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1127), .B(G330), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n319), .A2(new_n858), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n332), .B(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1135), .B1(new_n885), .B2(G330), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n903), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n885), .A2(G330), .A3(new_n1135), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n903), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1030), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n729), .B1(new_n201), .B2(new_n831), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n769), .A2(new_n202), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT117), .ZN(new_n1147));
  INV_X1    g0947(.A(G41), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n1148), .A3(new_n821), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1012), .B1(new_n229), .B2(new_n761), .C1(new_n224), .C2(new_n766), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n752), .A2(new_n426), .B1(new_n771), .B2(new_n770), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n756), .A2(new_n593), .B1(new_n750), .B2(new_n219), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n821), .A2(new_n1148), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G50), .B1(new_n259), .B2(new_n1148), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  MUX2_X1   g0956(.A(new_n1153), .B(new_n1156), .S(KEYINPUT58), .Z(new_n1157));
  OAI22_X1  g0957(.A1(new_n756), .A2(new_n1116), .B1(new_n750), .B2(new_n818), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1048), .A2(G137), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n1105), .B2(new_n766), .C1(new_n765), .C2(new_n1115), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G150), .C2(new_n781), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n926), .A2(G159), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n933), .C2(G124), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1157), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1145), .B1(new_n810), .B2(new_n1169), .C1(new_n1135), .C2(new_n742), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1126), .B1(new_n1144), .B2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1140), .A2(new_n1142), .A3(new_n1141), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1142), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n973), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(KEYINPUT118), .A3(new_n1170), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1093), .B1(new_n1095), .B2(new_n1089), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(KEYINPUT57), .A3(new_n1178), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n663), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1184), .ZN(G375));
  NAND2_X1  g0985(.A1(new_n1080), .A2(new_n1093), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n949), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1095), .A2(new_n1092), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n898), .A2(new_n741), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n729), .B1(new_n229), .B2(new_n831), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT119), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1147), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n779), .A2(G137), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n818), .B2(new_n756), .C1(new_n750), .C2(new_n1115), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n737), .B1(new_n1105), .B2(new_n771), .C1(new_n783), .C2(new_n765), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n752), .A2(new_n311), .B1(new_n761), .B2(new_n201), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n765), .A2(new_n219), .B1(new_n771), .B2(new_n763), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT120), .Z(new_n1201));
  OAI211_X1 g1001(.A(new_n1015), .B(new_n265), .C1(new_n217), .C2(new_n769), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n593), .A2(new_n750), .B1(new_n766), .B2(new_n770), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n756), .A2(new_n759), .B1(new_n752), .B2(new_n224), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1197), .A2(new_n1199), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1192), .B1(new_n810), .B2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  NAND2_X1  g1008(.A1(new_n1190), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1095), .B2(new_n1030), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1189), .A2(new_n1211), .ZN(G381));
  AOI21_X1  g1012(.A(G378), .B1(G375), .B2(KEYINPUT123), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(KEYINPUT123), .B2(G375), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1029), .A2(new_n1032), .A3(new_n794), .ZN(new_n1215));
  OR4_X1    g1015(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1215), .ZN(new_n1216));
  OR3_X1    g1016(.A1(new_n1214), .A2(G381), .A3(new_n1216), .ZN(G407));
  OAI211_X1 g1017(.A(G407), .B(G213), .C1(G343), .C2(new_n1214), .ZN(G409));
  NAND3_X1  g1018(.A1(new_n1177), .A2(new_n1184), .A3(G378), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1144), .A2(new_n1171), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1182), .A2(new_n1187), .A3(new_n1178), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(G378), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1219), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G213), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(G343), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1092), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1229), .A2(new_n663), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1092), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1188), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1233), .B2(new_n1211), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n835), .B(new_n1210), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1225), .A2(new_n1228), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT62), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT61), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1229), .A2(new_n663), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1188), .B2(new_n1231), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n835), .B1(new_n1241), .B2(new_n1210), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1233), .A2(G384), .A3(new_n1211), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1227), .A2(G2897), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1244), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G378), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n664), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1183), .A2(new_n1249), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1250), .B2(G378), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1245), .B(new_n1247), .C1(new_n1251), .C2(new_n1227), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1227), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1236), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1238), .A2(new_n1239), .A3(new_n1252), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n794), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1215), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n991), .A2(new_n992), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n972), .B2(new_n973), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1261), .A2(new_n948), .A3(G390), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n1261), .B2(new_n948), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1259), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(G390), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G387), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1215), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n1257), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n948), .A3(G390), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1264), .A2(new_n1270), .A3(KEYINPUT125), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT125), .B1(new_n1264), .B2(new_n1270), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1262), .A2(new_n1263), .A3(new_n1259), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1268), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1264), .A2(new_n1270), .A3(KEYINPUT125), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT126), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1274), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1256), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT124), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1237), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1247), .A2(new_n1245), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1239), .B(new_n1286), .C1(new_n1253), .C2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1237), .A2(new_n1283), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1282), .A2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(G375), .A2(new_n1223), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1219), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1236), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT127), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1294), .A2(new_n1296), .A3(new_n1219), .A4(new_n1236), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1301), .B(new_n1302), .ZN(G402));
endmodule


