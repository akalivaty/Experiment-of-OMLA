//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT68), .Z(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT67), .B(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT64), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n202), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(new_n221), .B2(new_n220), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n206), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n219), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT69), .B(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT5), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(G45), .C1(new_n255), .C2(KEYINPUT5), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT83), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(G41), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(KEYINPUT83), .A3(new_n254), .A4(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n251), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT76), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT76), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G257), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G264), .B2(new_n270), .ZN(new_n272));
  INV_X1    g0072(.A(G303), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n268), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n261), .A2(G270), .B1(new_n275), .B2(new_n251), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n256), .A2(new_n257), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n253), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n277), .A2(new_n260), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT84), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT84), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n258), .A2(new_n285), .A3(new_n281), .A4(new_n260), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT81), .B1(new_n262), .B2(G1), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT81), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n254), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G116), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n225), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT86), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n298), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n296), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT86), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(G116), .A4(new_n293), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G283), .ZN(new_n306));
  INV_X1    g0106(.A(G97), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n306), .B(new_n226), .C1(G33), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G116), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n296), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n308), .A2(KEYINPUT20), .A3(new_n296), .A4(new_n310), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n309), .B2(new_n301), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n305), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT79), .B(G190), .Z(new_n318));
  OAI211_X1 g0118(.A(new_n289), .B(new_n317), .C1(new_n288), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n305), .B2(new_n315), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT21), .B1(new_n321), .B2(new_n288), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n288), .A3(KEYINPUT21), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n316), .A2(G179), .A3(new_n287), .A4(new_n276), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n319), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT87), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n322), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT87), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n330), .A3(new_n319), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n281), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n279), .A2(new_n280), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n333), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G222), .A2(G1698), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n270), .A2(G223), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n274), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n265), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n267), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n336), .B1(new_n344), .B2(new_n213), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(G169), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n226), .A2(G33), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G20), .A2(G33), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n296), .A2(KEYINPUT70), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n295), .A2(new_n360), .A3(new_n225), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n358), .A2(new_n362), .B1(new_n202), .B2(new_n301), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n301), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n254), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G50), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT72), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n349), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n346), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(G190), .B2(new_n346), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n369), .A2(KEYINPUT9), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT9), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n363), .B2(new_n368), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n373), .C1(new_n374), .C2(new_n376), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n370), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n356), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n213), .B2(new_n353), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n362), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT75), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT11), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n384), .A2(KEYINPUT75), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n301), .A2(new_n210), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT12), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n302), .A2(G68), .A3(new_n365), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n338), .A2(new_n270), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n235), .A2(G1698), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n274), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n262), .B2(new_n307), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n251), .A2(new_n334), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(new_n251), .B1(G238), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n335), .B(KEYINPUT74), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n396), .B(G169), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT13), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(new_n405), .A3(G179), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n405), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n396), .B1(new_n413), .B2(G169), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n395), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(G200), .ZN(new_n416));
  INV_X1    g0216(.A(G190), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n394), .C1(new_n417), .C2(new_n413), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n335), .B1(new_n337), .B2(new_n212), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n274), .A2(G232), .A3(new_n270), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n274), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n420), .B1(new_n424), .B2(new_n251), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G169), .ZN(new_n426));
  INV_X1    g0226(.A(new_n350), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n356), .B1(G20), .B2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n354), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n297), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n302), .A2(G77), .A3(new_n365), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G77), .B2(new_n298), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OR3_X1    g0235(.A1(new_n426), .A2(new_n435), .A3(KEYINPUT73), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(new_n348), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT73), .B1(new_n426), .B2(new_n435), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n425), .A2(G190), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n435), .C1(new_n371), .C2(new_n425), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n381), .A2(new_n419), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n352), .A2(new_n365), .ZN(new_n443));
  INV_X1    g0243(.A(new_n352), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n443), .A2(new_n364), .B1(new_n301), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT77), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT7), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n268), .A2(new_n448), .A3(new_n226), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G68), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n268), .B2(new_n226), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT7), .B1(new_n453), .B2(G20), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT77), .A3(G68), .A4(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G58), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n210), .ZN(new_n458));
  OAI21_X1  g0258(.A(G20), .B1(new_n458), .B2(new_n201), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n356), .A2(G159), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(KEYINPUT16), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n448), .B1(new_n274), .B2(G20), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n461), .B1(new_n466), .B2(G68), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n296), .B1(new_n467), .B2(KEYINPUT16), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n446), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G223), .A2(G1698), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n338), .B2(G1698), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(new_n267), .A3(new_n263), .A4(new_n266), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G87), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n336), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n335), .B1(new_n235), .B2(new_n337), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n475), .A2(G179), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n338), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G223), .B2(G1698), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n474), .B1(new_n268), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n251), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n401), .A2(G232), .B1(new_n281), .B2(new_n334), .ZN(new_n482));
  AOI21_X1  g0282(.A(G169), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT78), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n482), .A3(new_n348), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(G169), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT18), .B1(new_n470), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n371), .B1(new_n481), .B2(new_n482), .ZN(new_n491));
  INV_X1    g0291(.A(new_n318), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT16), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n494), .B(new_n461), .C1(new_n452), .C2(new_n455), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n445), .B(new_n493), .C1(new_n495), .C2(new_n468), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n470), .A2(KEYINPUT17), .A3(new_n493), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n484), .A2(new_n488), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT18), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n461), .B1(new_n452), .B2(new_n455), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n468), .B1(new_n502), .B2(KEYINPUT16), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(new_n446), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n490), .A2(new_n498), .A3(new_n499), .A4(new_n504), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n442), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  INV_X1    g0308(.A(G244), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G1698), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(G238), .B2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n508), .B1(new_n268), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n251), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n254), .A2(new_n278), .A3(G45), .ZN(new_n514));
  INV_X1    g0314(.A(G45), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G1), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n336), .B(new_n514), .C1(G250), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G200), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n226), .B1(new_n262), .B2(new_n307), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n307), .A3(new_n423), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n353), .A2(KEYINPUT19), .A3(new_n307), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n263), .A2(new_n266), .A3(new_n226), .A4(new_n267), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n210), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(new_n296), .B1(new_n301), .B2(new_n429), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n359), .A2(new_n293), .A3(new_n298), .A4(new_n361), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G87), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n513), .A2(G190), .A3(new_n517), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n519), .A2(new_n528), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n296), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n430), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n429), .A2(new_n301), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n518), .A2(new_n320), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n513), .A2(new_n348), .A3(new_n517), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(KEYINPUT4), .A2(G244), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n267), .A2(new_n343), .A3(new_n542), .A4(new_n270), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT82), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n274), .A2(new_n545), .A3(new_n270), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n509), .A2(G1698), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n263), .A2(new_n266), .A3(new_n267), .A4(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n267), .A2(new_n343), .A3(G250), .A4(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n306), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n547), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n251), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n284), .A2(new_n286), .B1(new_n261), .B2(G257), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n348), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT7), .B1(new_n344), .B2(new_n226), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n448), .B(G20), .C1(new_n267), .C2(new_n343), .ZN(new_n561));
  OAI21_X1  g0361(.A(G107), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT80), .B(G107), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n307), .A2(new_n423), .A3(KEYINPUT6), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(KEYINPUT6), .B2(new_n307), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n563), .B(new_n565), .C1(KEYINPUT6), .C2(new_n307), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n356), .A2(G77), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n296), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n298), .A2(G97), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n529), .B2(new_n307), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n559), .A2(new_n320), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT85), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n556), .A2(new_n557), .A3(G190), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n571), .B2(new_n296), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n371), .B1(new_n556), .B2(new_n557), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n559), .A2(G200), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT85), .A3(new_n580), .A4(new_n579), .ZN(new_n585));
  AOI221_X4 g0385(.A(new_n541), .B1(new_n558), .B2(new_n577), .C1(new_n583), .C2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n529), .A2(new_n423), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n298), .A2(G107), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT90), .B(KEYINPUT25), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT23), .B1(new_n226), .B2(G107), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n423), .A3(G20), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT22), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n226), .A2(G87), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n344), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n599), .A2(new_n522), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n526), .A2(new_n604), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n602), .A2(new_n605), .B1(KEYINPUT88), .B2(KEYINPUT24), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n453), .A2(new_n226), .A3(new_n603), .ZN(new_n607));
  NOR2_X1   g0407(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n601), .A4(new_n598), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n296), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT89), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n613), .A3(new_n296), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n592), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n261), .A2(G264), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT91), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n269), .A2(G1698), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G250), .B2(G1698), .ZN(new_n619));
  INV_X1    g0419(.A(G294), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n268), .A2(new_n619), .B1(new_n262), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n251), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT91), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n261), .A2(new_n623), .A3(G264), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n617), .A2(new_n287), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n371), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n287), .A2(new_n616), .A3(new_n622), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(G190), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n615), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n613), .B1(new_n610), .B2(new_n296), .ZN(new_n630));
  AOI211_X1 g0430(.A(KEYINPUT89), .B(new_n297), .C1(new_n606), .C2(new_n609), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n591), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n627), .A2(G169), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n625), .B2(new_n348), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n332), .A2(new_n507), .A3(new_n586), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n370), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n490), .A2(new_n504), .ZN(new_n639));
  INV_X1    g0439(.A(new_n439), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n418), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n415), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n498), .A2(new_n499), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n639), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n378), .A2(new_n380), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n638), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n540), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n635), .A2(new_n329), .B1(new_n615), .B2(new_n628), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n586), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n580), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n261), .A2(G257), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n287), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n553), .B1(new_n550), .B2(new_n549), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n336), .B1(new_n656), .B2(new_n547), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n320), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(new_n658), .A3(new_n558), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n541), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT26), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n541), .B1(new_n659), .B2(KEYINPUT92), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT92), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n577), .A2(new_n663), .A3(new_n558), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT26), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT93), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI211_X1 g0467(.A(KEYINPUT93), .B(KEYINPUT26), .C1(new_n662), .C2(new_n664), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n652), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n649), .B1(new_n506), .B2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n254), .A2(new_n226), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n317), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n329), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n332), .B2(new_n680), .ZN(new_n682));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT94), .B1(new_n615), .B2(new_n678), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n632), .A2(new_n686), .A3(new_n677), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n636), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n632), .A2(new_n634), .A3(new_n677), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n678), .B1(new_n328), .B2(new_n322), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n688), .A2(new_n693), .B1(new_n635), .B2(new_n677), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n692), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n229), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n523), .A2(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n224), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n698), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n659), .A2(new_n541), .A3(KEYINPUT26), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n662), .A2(new_n664), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n677), .B1(new_n652), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT95), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n652), .A2(new_n706), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT95), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT29), .B1(new_n669), .B2(new_n678), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n624), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n623), .B1(new_n261), .B2(G264), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n622), .A2(new_n513), .A3(new_n517), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n559), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n276), .A2(G179), .A3(new_n287), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n718), .A2(new_n719), .A3(new_n556), .A4(new_n557), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n722), .ZN(new_n727));
  AOI21_X1  g0527(.A(G179), .B1(new_n513), .B2(new_n517), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n625), .A2(new_n559), .A3(new_n288), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n677), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n332), .A2(new_n636), .A3(new_n586), .A4(new_n678), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n715), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n703), .B1(new_n738), .B2(G1), .ZN(G364));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n684), .B(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n226), .A2(G13), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n254), .B1(new_n742), .B2(G45), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n698), .A2(KEYINPUT97), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT97), .ZN(new_n745));
  INV_X1    g0545(.A(new_n743), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n697), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n682), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(G330), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n741), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n748), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n274), .A2(new_n229), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n229), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n453), .A2(new_n696), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n224), .B2(new_n515), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n246), .A2(G45), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n225), .B1(G20), .B2(new_n320), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT98), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT98), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n752), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT99), .Z(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n417), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n226), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n774), .A2(new_n775), .B1(new_n620), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n772), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n318), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(G326), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT102), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n226), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n773), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n274), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n783), .A2(new_n417), .A3(G200), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n786), .B1(new_n787), .B2(new_n788), .C1(new_n273), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n772), .A2(new_n371), .A3(new_n492), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G322), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT101), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n779), .B2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n779), .A2(new_n794), .A3(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  OAI21_X1  g0599(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(new_n210), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n274), .B1(new_n423), .B2(new_n788), .C1(new_n791), .C2(new_n457), .ZN(new_n802));
  INV_X1    g0602(.A(new_n774), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G77), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n780), .A2(G50), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n784), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT100), .B(KEYINPUT32), .Z(new_n808));
  XNOR2_X1  g0608(.A(new_n807), .B(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n777), .A2(new_n307), .B1(new_n789), .B2(new_n522), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n804), .A2(new_n805), .A3(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n782), .A2(new_n800), .B1(new_n801), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n770), .B1(new_n813), .B2(new_n764), .ZN(new_n814));
  INV_X1    g0614(.A(new_n767), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n749), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n751), .A2(new_n816), .ZN(G396));
  INV_X1    g0617(.A(KEYINPUT103), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n439), .A2(new_n818), .A3(new_n441), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n677), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n669), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n677), .B1(new_n432), .B2(new_n434), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(KEYINPUT103), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n439), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n669), .B2(new_n678), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n748), .B1(new_n829), .B2(new_n736), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(KEYINPUT104), .B1(new_n736), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT104), .B2(new_n830), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n792), .A2(G143), .B1(new_n803), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(new_n780), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n833), .B1(new_n834), .B2(new_n835), .C1(new_n798), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n453), .B1(new_n839), .B2(new_n784), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n788), .A2(new_n210), .ZN(new_n841));
  INV_X1    g0641(.A(new_n777), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(G58), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n202), .B2(new_n789), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n838), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n798), .A2(new_n787), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n344), .B1(new_n784), .B2(new_n775), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n522), .A2(new_n788), .B1(new_n789), .B2(new_n423), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(G97), .C2(new_n842), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n309), .B2(new_n774), .C1(new_n620), .C2(new_n791), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n846), .B(new_n850), .C1(G303), .C2(new_n780), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n764), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n764), .A2(new_n765), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n748), .B1(new_n853), .B2(new_n213), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n854), .C1(new_n766), .C2(new_n827), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n832), .A2(new_n855), .ZN(G384));
  OAI211_X1 g0656(.A(new_n224), .B(G77), .C1(new_n457), .C2(new_n210), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n202), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n254), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n567), .A2(new_n568), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT35), .ZN(new_n861));
  OAI211_X1 g0661(.A(G116), .B(new_n227), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT36), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n500), .B1(new_n503), .B2(new_n446), .ZN(new_n867));
  INV_X1    g0667(.A(new_n675), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n503), .B2(new_n446), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n869), .A3(new_n496), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n362), .B1(new_n502), .B2(KEYINPUT16), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT105), .B(new_n362), .C1(new_n502), .C2(KEYINPUT16), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n463), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n445), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n868), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n500), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n496), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n871), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n675), .B1(new_n876), .B2(new_n445), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n505), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n866), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n883), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  INV_X1    g0686(.A(new_n496), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n877), .B2(new_n500), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n878), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n885), .C1(new_n889), .C2(new_n871), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n495), .B1(new_n872), .B2(new_n873), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n446), .B1(new_n893), .B2(new_n875), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n496), .B1(new_n894), .B2(new_n489), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  INV_X1    g0696(.A(new_n871), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n866), .B(new_n883), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n870), .B(KEYINPUT37), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n505), .B(new_n868), .C1(new_n446), .C2(new_n503), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n892), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n415), .A2(new_n677), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n891), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n868), .B1(new_n490), .B2(new_n504), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n884), .A2(new_n890), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n439), .A2(new_n677), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n669), .B2(new_n820), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n415), .A2(new_n418), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n395), .A3(new_n677), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n415), .B(new_n418), .C1(new_n394), .C2(new_n678), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n906), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n905), .A2(new_n916), .A3(KEYINPUT106), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT106), .B1(new_n905), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n648), .B1(new_n714), .B2(new_n507), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT107), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n883), .B1(new_n896), .B2(new_n897), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n901), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n826), .B1(new_n911), .B2(new_n912), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n735), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT40), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n735), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n896), .A2(new_n897), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n931), .B2(new_n885), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n930), .B1(new_n932), .B2(new_n898), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n934), .A2(new_n507), .A3(new_n735), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n507), .B2(new_n735), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n935), .A2(new_n936), .A3(new_n683), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n922), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT108), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n939), .B1(new_n254), .B2(new_n742), .C1(new_n922), .C2(new_n937), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(KEYINPUT108), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n865), .B1(new_n940), .B2(new_n941), .ZN(G367));
  INV_X1    g0742(.A(new_n789), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT46), .B1(new_n943), .B2(G116), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(KEYINPUT46), .A3(G116), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n791), .B2(new_n273), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n944), .B(new_n946), .C1(G283), .C2(new_n803), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n453), .B1(G317), .B2(new_n785), .ZN(new_n948));
  INV_X1    g0748(.A(new_n788), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(G97), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(new_n423), .C2(new_n777), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G311), .B2(new_n780), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n947), .B(new_n952), .C1(new_n620), .C2(new_n798), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n798), .A2(new_n806), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n791), .A2(new_n836), .B1(new_n210), .B2(new_n777), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT112), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n780), .A2(G143), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n788), .A2(new_n213), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n274), .B1(new_n784), .B2(new_n834), .C1(new_n457), .C2(new_n789), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(new_n803), .C2(G50), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n953), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT47), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n764), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n528), .A2(new_n531), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n677), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n540), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n533), .A2(new_n540), .A3(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n767), .A3(new_n970), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n768), .B1(new_n229), .B2(new_n429), .C1(new_n241), .C2(new_n757), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT111), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n974), .A2(new_n975), .A3(new_n748), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n966), .A2(new_n971), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n688), .A2(new_n693), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n688), .A2(new_n689), .A3(new_n693), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(KEYINPUT110), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(KEYINPUT110), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n741), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n684), .B2(new_n982), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n583), .A2(new_n585), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n985), .B(new_n659), .C1(new_n580), .C2(new_n678), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n577), .A2(new_n558), .A3(new_n677), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n694), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n694), .A2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(KEYINPUT109), .A3(new_n692), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n692), .A2(KEYINPUT109), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n990), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n984), .A2(new_n995), .A3(new_n738), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(new_n738), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n697), .B(KEYINPUT41), .Z(new_n1000));
  OAI21_X1  g0800(.A(new_n743), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n986), .A2(new_n635), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n677), .B1(new_n1002), .B2(new_n659), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n979), .A2(new_n988), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(KEYINPUT42), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT42), .B2(new_n1004), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n969), .A2(new_n970), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1006), .A2(KEYINPUT43), .A3(new_n1007), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n691), .A2(new_n988), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1013), .B(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n978), .B1(new_n1001), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n982), .A2(new_n684), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1019), .B(new_n746), .C1(new_n741), .C2(new_n982), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n753), .A2(new_n699), .B1(G107), .B2(new_n229), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n238), .A2(new_n515), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n699), .ZN(new_n1023));
  AOI211_X1 g0823(.A(G45), .B(new_n1023), .C1(G68), .C2(G77), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n350), .A2(G50), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n757), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1021), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n752), .B1(new_n1028), .B2(new_n769), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n453), .B1(new_n836), .B2(new_n784), .C1(new_n774), .C2(new_n210), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G50), .B2(new_n792), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n950), .B1(new_n213), .B2(new_n789), .C1(new_n429), .C2(new_n777), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n780), .B2(G159), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(new_n444), .C2(new_n798), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n453), .B1(G326), .B2(new_n785), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n777), .A2(new_n787), .B1(new_n789), .B2(new_n620), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n792), .A2(G317), .B1(new_n803), .B2(G303), .ZN(new_n1037));
  INV_X1    g0837(.A(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n835), .C1(new_n798), .C2(new_n775), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1035), .B1(new_n309), .B2(new_n788), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1029), .B1(new_n1046), .B2(new_n764), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n690), .B2(new_n815), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1020), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n984), .A2(new_n738), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1019), .B1(new_n741), .B2(new_n982), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n697), .B1(new_n1051), .B2(new_n737), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1049), .B1(new_n1050), .B2(new_n1052), .ZN(G393));
  NOR2_X1   g0853(.A1(new_n994), .A2(new_n692), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n691), .B1(new_n990), .B2(new_n993), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1054), .A2(new_n1055), .B1(new_n1051), .B2(new_n737), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n998), .A2(new_n1056), .A3(new_n697), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT116), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT116), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n998), .A2(new_n1056), .A3(new_n1059), .A4(new_n697), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n249), .A2(new_n756), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n768), .B1(new_n307), .B2(new_n229), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n798), .A2(new_n202), .B1(new_n350), .B2(new_n774), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT114), .Z(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n780), .B1(new_n792), .B2(G159), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n777), .A2(new_n213), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G87), .B2(new_n949), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n268), .B1(new_n785), .B2(G143), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n210), .C2(new_n789), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G317), .A2(new_n780), .B1(new_n792), .B2(G311), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT52), .Z(new_n1074));
  NOR2_X1   g0874(.A1(new_n798), .A2(new_n273), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n274), .B1(new_n949), .B2(G107), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n309), .B2(new_n777), .C1(new_n774), .C2(new_n620), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n789), .A2(new_n787), .B1(new_n784), .B2(new_n1038), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT115), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1075), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1065), .A2(new_n1072), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n764), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n752), .B1(new_n1062), .B2(new_n1063), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n767), .B2(new_n988), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT113), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n743), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR3_X1    g0887(.A1(new_n1054), .A2(new_n1086), .A3(new_n1055), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1061), .A2(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(new_n901), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n890), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n908), .B1(new_n707), .B2(new_n827), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n903), .C1(new_n914), .C2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n903), .B1(new_n909), .B2(new_n914), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT117), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(KEYINPUT117), .B(new_n903), .C1(new_n909), .C2(new_n914), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n890), .B2(new_n1091), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n932), .A2(new_n898), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(KEYINPUT39), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1094), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n683), .B1(new_n733), .B2(new_n734), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n827), .A3(new_n913), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n891), .A2(new_n902), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(new_n1106), .A3(new_n1094), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n765), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n791), .A2(new_n309), .B1(new_n774), .B2(new_n307), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n344), .B1(new_n784), .B2(new_n620), .C1(new_n522), .C2(new_n789), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1114), .A2(new_n841), .A3(new_n1068), .A4(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n787), .B2(new_n835), .C1(new_n798), .C2(new_n423), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT120), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n344), .B1(new_n785), .B2(G125), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n202), .B2(new_n788), .C1(new_n806), .C2(new_n777), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G128), .B2(new_n780), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n791), .A2(new_n839), .B1(new_n774), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n789), .A2(new_n836), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1126));
  XNOR2_X1  g0926(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1122), .B(new_n1128), .C1(new_n834), .C2(new_n798), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1119), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1131), .A2(new_n764), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n748), .B(new_n1132), .C1(new_n444), .C2(new_n853), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1112), .A2(new_n746), .B1(new_n1113), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n506), .A2(new_n736), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n920), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1104), .A2(new_n827), .A3(new_n913), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n913), .B1(new_n1104), .B2(new_n827), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1138), .A2(new_n1139), .B1(new_n821), .B2(new_n908), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n914), .B1(new_n736), .B2(new_n826), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1105), .A3(new_n1093), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n697), .B1(new_n1112), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n648), .B(new_n1135), .C1(new_n714), .C2(new_n507), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1134), .B1(new_n1145), .B2(new_n1149), .ZN(G378));
  NAND2_X1  g0950(.A1(new_n369), .A2(new_n868), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT55), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1151), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT123), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n381), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n381), .A2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1154), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1154), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1156), .A3(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(new_n766), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n748), .B1(new_n853), .B2(new_n202), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n777), .A2(new_n836), .B1(new_n789), .B2(new_n1123), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n792), .A2(G128), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G137), .C2(new_n803), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n780), .A2(G125), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n839), .C2(new_n798), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n949), .A2(G159), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n268), .A2(new_n255), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n774), .A2(new_n429), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G107), .C2(new_n792), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n777), .A2(new_n210), .B1(new_n787), .B2(new_n784), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n949), .A2(G58), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n213), .B2(new_n789), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G116), .C2(new_n780), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1178), .B(new_n1182), .C1(new_n307), .C2(new_n798), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1176), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT121), .Z(new_n1188));
  AND4_X1   g0988(.A1(new_n1175), .A2(new_n1185), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1165), .B1(new_n1189), .B2(new_n1082), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1164), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1163), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n934), .B2(G330), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n683), .B(new_n1163), .C1(new_n927), .C2(new_n933), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n918), .A2(new_n917), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n905), .A2(new_n916), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT106), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n926), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n928), .B1(new_n1092), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n929), .B1(new_n884), .B2(new_n890), .ZN(new_n1201));
  OAI21_X1  g1001(.A(G330), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1163), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n905), .A2(new_n916), .A3(KEYINPUT106), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n934), .A2(G330), .A3(new_n1192), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1198), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1195), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1191), .B1(new_n1207), .B2(new_n746), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1110), .A2(new_n1106), .A3(new_n1094), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1106), .B1(new_n1110), .B2(new_n1094), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1144), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1212), .A2(new_n1146), .B1(new_n1195), .B2(new_n1206), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n698), .B1(new_n1213), .B2(KEYINPUT57), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1146), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1207), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT57), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1209), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1000), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1148), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1147), .A2(new_n746), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n748), .B1(new_n853), .B2(new_n210), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT124), .Z(new_n1226));
  OAI22_X1  g1026(.A1(new_n791), .A2(new_n787), .B1(new_n774), .B2(new_n423), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n344), .B1(new_n784), .B2(new_n273), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n777), .A2(new_n429), .B1(new_n789), .B2(new_n307), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1227), .A2(new_n958), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n620), .B2(new_n835), .C1(new_n309), .C2(new_n798), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1180), .B1(new_n806), .B2(new_n789), .C1(new_n202), .C2(new_n777), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n780), .B2(G132), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n268), .B1(new_n785), .B2(G128), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n774), .B2(new_n836), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G137), .B2(new_n792), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(new_n798), .C2(new_n1123), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1231), .A2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1226), .B1(new_n1082), .B2(new_n1238), .C1(new_n913), .C2(new_n766), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1224), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1223), .A2(new_n1241), .ZN(G381));
  INV_X1    g1042(.A(G378), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1219), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G396), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1049), .B(new_n1245), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1246), .A2(G381), .A3(G384), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G387), .A2(new_n1244), .A3(G390), .A4(new_n1247), .ZN(G407));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n697), .B1(new_n1221), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1253), .A2(new_n1144), .A3(KEYINPUT125), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1250), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n1148), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1252), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G384), .A3(new_n1241), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT125), .B1(new_n1253), .B2(new_n1144), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(new_n1255), .A3(new_n1148), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1251), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1263), .B2(new_n1240), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1266), .A2(G2897), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1259), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1207), .B(KEYINPUT57), .C1(new_n1137), .C2(new_n1149), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n697), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1207), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1208), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1208), .B1(new_n1216), .B2(new_n1000), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1243), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1266), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1270), .B1(new_n1277), .B2(KEYINPUT126), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1213), .A2(new_n1222), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G378), .B1(new_n1208), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1219), .B2(G378), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(new_n1282), .B2(new_n1266), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1246), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1061), .A2(new_n1286), .A3(new_n1089), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1061), .B2(new_n1089), .ZN(new_n1288));
  OAI21_X1  g1088(.A(G387), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G390), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1061), .A2(new_n1286), .A3(new_n1089), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1017), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1289), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1266), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1259), .A2(new_n1264), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1295), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1298), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1284), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1277), .A2(new_n1304), .A3(new_n1298), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1294), .B1(new_n1277), .B2(new_n1270), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1277), .B2(new_n1298), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1303), .B1(new_n1308), .B2(new_n1310), .ZN(G405));
  NOR2_X1   g1111(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1312));
  OR2_X1    g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1274), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1219), .A2(G378), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1313), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1313), .B2(new_n1318), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G402));
endmodule


