//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT66), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n213), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT7), .B1(new_n252), .B2(new_n214), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  AOI211_X1 g0054(.A(new_n254), .B(G20), .C1(new_n249), .C2(new_n251), .ZN(new_n255));
  OAI21_X1  g0055(.A(G68), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  INV_X1    g0057(.A(G68), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n259), .B2(new_n201), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G159), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT16), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n247), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT70), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n254), .B1(new_n269), .B2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n263), .B1(new_n272), .B2(G68), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n268), .B1(new_n273), .B2(KEYINPUT16), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n275));
  NOR4_X1   g0075(.A1(new_n275), .A2(new_n263), .A3(KEYINPUT70), .A4(new_n266), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n267), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT8), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n213), .A3(new_n245), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n284), .A2(new_n286), .B1(new_n285), .B2(new_n281), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n293), .A3(G274), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n282), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(G232), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(G226), .A2(G1698), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n249), .A2(new_n251), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G87), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n249), .A2(new_n251), .A3(G223), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT71), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n249), .A2(new_n251), .A3(new_n298), .A4(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n300), .A2(new_n301), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G200), .B2(new_n308), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n277), .A2(new_n288), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT17), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n277), .A2(KEYINPUT17), .A3(new_n288), .A4(new_n311), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT74), .B1(new_n314), .B2(new_n315), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n285), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n258), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n258), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n214), .A2(G33), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n218), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT11), .A3(new_n246), .ZN(new_n325));
  INV_X1    g0125(.A(new_n286), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G68), .A3(new_n283), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT11), .B1(new_n324), .B2(new_n246), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n249), .A2(new_n251), .A3(G232), .A4(G1698), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n249), .A2(new_n251), .A3(G226), .A4(new_n302), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G97), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n336), .A2(new_n307), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT68), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n291), .A2(new_n293), .A3(new_n339), .A4(G274), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n293), .A2(G238), .A3(new_n295), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n337), .A2(new_n342), .A3(KEYINPUT13), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n341), .ZN(new_n345));
  INV_X1    g0145(.A(G274), .ZN(new_n346));
  INV_X1    g0146(.A(new_n213), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n292), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n339), .B1(new_n348), .B2(new_n291), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n336), .A2(new_n307), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n332), .B(G169), .C1(new_n343), .C2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT13), .B1(new_n337), .B2(new_n342), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n344), .A3(new_n351), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G179), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n355), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n332), .B1(new_n358), .B2(G169), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n331), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n269), .A2(G222), .A3(new_n302), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n269), .A2(G223), .A3(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n218), .C2(new_n269), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n307), .ZN(new_n364));
  INV_X1    g0164(.A(new_n294), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n307), .A2(new_n291), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(G226), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n323), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n281), .A2(new_n371), .B1(G150), .B2(new_n261), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n203), .A2(G20), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n247), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n283), .A2(G50), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n286), .A2(new_n375), .B1(G50), .B2(new_n285), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n368), .A2(G179), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(KEYINPUT9), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT9), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n374), .B2(new_n376), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n364), .A2(G190), .A3(new_n367), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n368), .A2(G200), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n388), .A2(new_n387), .A3(new_n384), .A4(new_n382), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n381), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n354), .A2(G190), .A3(new_n355), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT69), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n358), .B2(G200), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  AOI211_X1 g0196(.A(KEYINPUT69), .B(new_n396), .C1(new_n354), .C2(new_n355), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n330), .B(new_n393), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(KEYINPUT8), .B(G58), .ZN(new_n399));
  INV_X1    g0199(.A(new_n261), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(new_n214), .B2(new_n218), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n323), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n246), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT67), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n218), .B1(new_n282), .B2(G20), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n326), .A2(new_n406), .B1(new_n218), .B2(new_n319), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n269), .A2(G232), .A3(new_n302), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n269), .A2(G238), .A3(G1698), .ZN(new_n410));
  INV_X1    g0210(.A(G107), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n269), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n307), .ZN(new_n413));
  INV_X1    g0213(.A(new_n217), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n365), .B1(new_n414), .B2(new_n366), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n369), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n408), .B(new_n417), .C1(G179), .C2(new_n416), .ZN(new_n418));
  INV_X1    g0218(.A(new_n416), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G190), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(G200), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n405), .A4(new_n407), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AND4_X1   g0223(.A1(new_n360), .A2(new_n392), .A3(new_n398), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n256), .A2(KEYINPUT16), .A3(new_n264), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT70), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n273), .A2(new_n268), .A3(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n287), .B1(new_n428), .B2(new_n267), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n306), .A2(new_n307), .ZN(new_n431));
  INV_X1    g0231(.A(new_n297), .ZN(new_n432));
  AOI21_X1  g0232(.A(G169), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(G179), .B(new_n297), .C1(new_n306), .C2(new_n307), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT72), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G179), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(G169), .C2(new_n308), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT73), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n435), .B2(new_n439), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n430), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT18), .B(new_n430), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n318), .A2(new_n424), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n249), .A2(new_n251), .A3(G264), .A4(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n249), .A2(new_n251), .A3(G257), .A4(new_n302), .ZN(new_n450));
  INV_X1    g0250(.A(G303), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(new_n450), .C1(new_n451), .C2(new_n269), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n452), .A2(new_n307), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n290), .A2(G1), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n348), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n293), .ZN(new_n460));
  INV_X1    g0260(.A(G270), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT80), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n452), .A2(new_n307), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n307), .B1(new_n454), .B2(new_n455), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G270), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n456), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n285), .A2(G116), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT75), .B1(new_n248), .B2(G1), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT75), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n282), .A3(G33), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n286), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n469), .B1(new_n474), .B2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n214), .C1(G33), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G20), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n246), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n478), .A2(new_n246), .A3(KEYINPUT20), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n369), .B1(new_n475), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n463), .A2(new_n468), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n453), .A2(new_n436), .A3(new_n462), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n475), .A2(new_n485), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n463), .A2(new_n486), .A3(KEYINPUT21), .A4(new_n468), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n463), .A2(new_n468), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n491), .B1(new_n495), .B2(G190), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n396), .B2(new_n495), .ZN(new_n497));
  XNOR2_X1  g0297(.A(G97), .B(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n477), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n411), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n272), .A2(G107), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(G97), .B1(new_n473), .B2(new_n286), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n285), .A2(new_n477), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT76), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(KEYINPUT76), .A3(new_n508), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n506), .A2(new_n246), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n249), .A2(new_n251), .A3(G244), .A4(new_n302), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT77), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n515), .A2(KEYINPUT4), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n269), .A2(G244), .A3(new_n516), .A4(new_n302), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n476), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n307), .ZN(new_n522));
  INV_X1    g0322(.A(G257), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n456), .B1(new_n460), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n521), .B2(new_n307), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G190), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n513), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n511), .A2(new_n512), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n498), .A2(new_n499), .B1(new_n411), .B2(new_n501), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n532), .A2(new_n214), .B1(new_n218), .B2(new_n400), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n411), .B1(new_n270), .B2(new_n271), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n246), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n526), .A2(new_n369), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n528), .A2(new_n436), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n269), .A2(new_n214), .A3(G68), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n323), .B2(new_n477), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n477), .A3(new_n411), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT79), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT79), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(new_n545), .A3(new_n477), .A4(new_n411), .ZN(new_n549));
  NAND3_X1  g0349(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(new_n549), .B1(new_n214), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n246), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n402), .A2(new_n319), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n474), .A2(G87), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n293), .A2(G274), .A3(new_n454), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  OR2_X1    g0358(.A1(G238), .A2(G1698), .ZN(new_n559));
  INV_X1    g0359(.A(G244), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n558), .B1(new_n562), .B2(new_n252), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n557), .B1(new_n563), .B2(new_n307), .ZN(new_n564));
  OAI21_X1  g0364(.A(G250), .B1(new_n290), .B2(G1), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT78), .B1(new_n307), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n565), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT78), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n293), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n564), .A2(G190), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n396), .B1(new_n564), .B2(new_n570), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n556), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n402), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n474), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n552), .A2(new_n553), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n564), .A2(G179), .A3(new_n570), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n369), .B1(new_n564), .B2(new_n570), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n494), .A2(new_n497), .A3(new_n540), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n285), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n411), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n474), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n249), .A2(new_n251), .A3(new_n214), .A4(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT22), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n269), .A2(new_n592), .A3(new_n214), .A4(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n558), .A2(G20), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n214), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n411), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT24), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n594), .A2(new_n602), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n589), .B1(new_n604), .B2(new_n246), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n249), .A2(new_n251), .A3(G257), .A4(G1698), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(new_n302), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G33), .A2(G294), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n307), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n466), .A2(G264), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n456), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n369), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G179), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n584), .B1(new_n605), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n594), .A2(new_n602), .A3(new_n599), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n602), .B1(new_n594), .B2(new_n599), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n246), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n588), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n612), .A2(G179), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n307), .A2(new_n609), .B1(new_n466), .B2(G264), .ZN(new_n621));
  AOI21_X1  g0421(.A(G169), .B1(new_n621), .B2(new_n456), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n623), .A3(KEYINPUT81), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(G190), .A3(new_n456), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n612), .A2(G200), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n618), .A2(new_n588), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n615), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT82), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n615), .A2(KEYINPUT82), .A3(new_n624), .A4(new_n627), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n583), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n448), .A2(new_n632), .ZN(G372));
  AND2_X1   g0433(.A1(new_n389), .A2(new_n391), .ZN(new_n634));
  INV_X1    g0434(.A(new_n317), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n393), .A2(new_n330), .ZN(new_n636));
  INV_X1    g0436(.A(new_n395), .ZN(new_n637));
  INV_X1    g0437(.A(new_n397), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n360), .B1(new_n639), .B2(new_n418), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n315), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n435), .A2(new_n439), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n429), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n644), .B(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n634), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n381), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n530), .A2(new_n539), .A3(new_n627), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n619), .A2(new_n623), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(new_n489), .A3(new_n492), .A4(new_n493), .ZN(new_n651));
  INV_X1    g0451(.A(new_n571), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n652), .A2(new_n555), .A3(new_n572), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT83), .B1(new_n578), .B2(new_n579), .ZN(new_n654));
  INV_X1    g0454(.A(new_n557), .ZN(new_n655));
  NOR2_X1   g0455(.A1(G238), .A2(G1698), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n560), .B2(G1698), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n269), .B1(G33), .B2(G116), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n293), .ZN(new_n659));
  INV_X1    g0459(.A(new_n570), .ZN(new_n660));
  OAI21_X1  g0460(.A(G169), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT83), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n564), .A2(G179), .A3(new_n570), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n653), .B1(new_n665), .B2(new_n577), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n649), .A2(new_n651), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT83), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n577), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .A4(new_n574), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n581), .B2(new_n539), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n448), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n648), .A2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G1), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n214), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G213), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(new_n491), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n494), .A2(new_n497), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(KEYINPUT86), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT86), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n494), .A2(new_n692), .A3(new_n497), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n494), .A2(new_n689), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT87), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(KEYINPUT87), .A3(new_n695), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n679), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n630), .A2(new_n631), .ZN(new_n701));
  INV_X1    g0501(.A(new_n688), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n605), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n650), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n688), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n494), .A2(new_n688), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n702), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(G399));
  NAND3_X1  g0512(.A1(new_n547), .A2(new_n479), .A3(new_n549), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n207), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(G1), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n211), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n721), .B(new_n702), .C1(new_n667), .C2(new_n675), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n493), .A2(new_n492), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n615), .A2(new_n723), .A3(new_n624), .A4(new_n489), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n666), .A3(new_n649), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n666), .A2(new_n671), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT26), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n581), .A2(new_n539), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(new_n672), .B1(new_n577), .B2(new_n665), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(new_n702), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n722), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AND4_X1   g0535(.A1(new_n611), .A2(new_n564), .A3(new_n610), .A4(new_n570), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n490), .A2(new_n736), .A3(new_n528), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n490), .A2(new_n736), .A3(KEYINPUT30), .A4(new_n528), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(G179), .B1(new_n564), .B2(new_n570), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n463), .A2(new_n468), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n612), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT90), .B1(new_n744), .B2(new_n528), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT90), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n526), .A2(new_n746), .A3(new_n612), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n688), .B(new_n735), .C1(new_n741), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n688), .B1(new_n741), .B2(new_n748), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n583), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n701), .A2(new_n754), .A3(new_n702), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n733), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n720), .B1(new_n759), .B2(G1), .ZN(G364));
  INV_X1    g0560(.A(new_n699), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT87), .B1(new_n694), .B2(new_n695), .ZN(new_n762));
  OAI21_X1  g0562(.A(G330), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n698), .A2(new_n679), .A3(new_n699), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n680), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n282), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n716), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n213), .B1(G20), .B2(new_n369), .ZN(new_n771));
  NAND2_X1  g0571(.A1(G20), .A2(G179), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT92), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n396), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n309), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n214), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n775), .A2(G326), .B1(G294), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n773), .A2(new_n309), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n779), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT94), .Z(new_n785));
  NOR2_X1   g0585(.A1(new_n214), .A2(G179), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n252), .B1(new_n787), .B2(new_n451), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT95), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n786), .A2(new_n309), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(new_n309), .A3(new_n396), .ZN(new_n792));
  INV_X1    g0592(.A(G329), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n774), .A2(G200), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(G322), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n781), .A2(new_n396), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(G317), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n796), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n785), .A2(new_n789), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n775), .ZN(new_n803));
  INV_X1    g0603(.A(new_n795), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n202), .A2(new_n803), .B1(new_n804), .B2(new_n257), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n258), .A2(new_n798), .B1(new_n783), .B2(new_n218), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n792), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  INV_X1    g0609(.A(new_n790), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n252), .B1(new_n810), .B2(G107), .ZN(new_n811));
  INV_X1    g0611(.A(new_n787), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n778), .A2(G97), .B1(new_n812), .B2(G87), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n805), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n771), .B1(new_n802), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n269), .A2(new_n207), .ZN(new_n818));
  INV_X1    g0618(.A(G355), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n818), .A2(new_n819), .B1(G116), .B2(new_n207), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n238), .A2(new_n290), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n715), .A2(new_n269), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n290), .B2(new_n212), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n820), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n771), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n768), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT91), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n817), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n696), .B2(new_n828), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n770), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  NOR2_X1   g0636(.A1(new_n771), .A2(new_n826), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n769), .B1(new_n218), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n418), .A2(new_n688), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n688), .A2(new_n408), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n422), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n418), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G294), .A2(new_n795), .B1(new_n775), .B2(G303), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n791), .B2(new_n798), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n783), .A2(new_n479), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n252), .B1(new_n792), .B2(new_n780), .C1(new_n777), .C2(new_n477), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n545), .A2(new_n790), .B1(new_n787), .B2(new_n411), .ZN(new_n847));
  NOR4_X1   g0647(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n795), .B1(new_n782), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n803), .C1(new_n851), .C2(new_n798), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT34), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n269), .B1(new_n792), .B2(new_n854), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n202), .A2(new_n787), .B1(new_n790), .B2(new_n258), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(G58), .C2(new_n778), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n848), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n771), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n838), .B1(new_n842), .B2(new_n827), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n757), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n842), .B1(new_n676), .B2(new_n702), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n702), .B(new_n842), .C1(new_n667), .C2(new_n675), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n769), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n866), .B1(new_n868), .B2(KEYINPUT97), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(KEYINPUT97), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(G384));
  INV_X1    g0672(.A(new_n645), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n644), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n686), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n267), .A2(KEYINPUT98), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n246), .B1(new_n273), .B2(KEYINPUT16), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT98), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n428), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n288), .ZN(new_n881));
  INV_X1    g0681(.A(new_n686), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n445), .A2(new_n446), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n635), .A2(new_n641), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(new_n435), .A3(new_n439), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n312), .A3(new_n883), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n312), .B1(new_n429), .B2(new_n686), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n889), .A2(KEYINPUT37), .B1(new_n891), .B2(new_n443), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n883), .B1(new_n318), .B2(new_n447), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n895), .A2(new_n896), .A3(new_n892), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n839), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n863), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n688), .A2(new_n331), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n360), .A2(new_n398), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n360), .B2(new_n398), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n875), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n890), .B2(new_n644), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT99), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n891), .A2(new_n443), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT99), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(KEYINPUT37), .C1(new_n890), .C2(new_n644), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT100), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT100), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n430), .A2(new_n882), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n314), .A2(new_n315), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n646), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(new_n917), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n896), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n318), .A2(new_n447), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n892), .B1(new_n925), .B2(new_n884), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT39), .B1(new_n926), .B2(KEYINPUT38), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n896), .B1(new_n895), .B2(new_n892), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n924), .A2(new_n927), .B1(new_n930), .B2(KEYINPUT39), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n357), .A2(new_n359), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n331), .A3(new_n702), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n908), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n721), .B1(new_n730), .B2(new_n702), .ZN(new_n935));
  INV_X1    g0735(.A(new_n722), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n448), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n648), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT101), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n934), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n752), .A2(new_n734), .ZN(new_n941));
  OAI211_X1 g0741(.A(KEYINPUT31), .B(new_n688), .C1(new_n741), .C2(new_n748), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n755), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n842), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n904), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n921), .B1(new_n914), .B2(new_n915), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT38), .B1(new_n949), .B2(new_n917), .ZN(new_n950));
  OAI211_X1 g0750(.A(KEYINPUT40), .B(new_n948), .C1(new_n950), .C2(new_n897), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n894), .B2(new_n897), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT40), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n318), .A2(new_n424), .A3(new_n447), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n941), .A2(new_n942), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n632), .B2(new_n702), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n955), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n956), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(G330), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n940), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(KEYINPUT102), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(KEYINPUT102), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n940), .A2(new_n962), .B1(new_n282), .B2(new_n765), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(G116), .A3(new_n215), .A4(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT36), .Z(new_n971));
  OR3_X1    g0771(.A1(new_n211), .A2(new_n218), .A3(new_n259), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n202), .A2(G68), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n282), .B(G13), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n967), .A2(new_n971), .A3(new_n974), .ZN(G367));
  INV_X1    g0775(.A(new_n666), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n702), .A2(new_n556), .ZN(new_n977));
  MUX2_X1   g0777(.A(new_n976), .B(new_n670), .S(new_n977), .Z(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n710), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n540), .B1(new_n513), .B2(new_n702), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n671), .A2(new_n688), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n615), .A2(new_n624), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n688), .B1(new_n988), .B2(new_n539), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n985), .B2(KEYINPUT42), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n980), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n978), .A2(new_n979), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n984), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n707), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n716), .B(KEYINPUT41), .Z(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT103), .B1(new_n706), .B2(new_n709), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n763), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n700), .A2(new_n998), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n981), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n981), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n759), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT104), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n710), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(KEYINPUT104), .A3(new_n759), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n710), .A2(new_n711), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1012), .A2(KEYINPUT44), .A3(new_n994), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT44), .B1(new_n1012), .B2(new_n994), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n994), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT45), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1012), .A2(new_n1017), .A3(new_n994), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n707), .B1(new_n1013), .B2(new_n1014), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1016), .A2(new_n1018), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1020), .A2(new_n700), .A3(new_n706), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1007), .A2(new_n1011), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n997), .B1(new_n1022), .B2(new_n759), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n996), .B1(new_n1023), .B2(new_n767), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n829), .B1(new_n207), .B2(new_n402), .C1(new_n234), .C2(new_n823), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n777), .A2(new_n258), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n269), .B1(new_n792), .B2(new_n850), .C1(new_n218), .C2(new_n790), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G58), .C2(new_n812), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n797), .A2(G159), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n775), .A2(G143), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G50), .A2(new_n782), .B1(new_n795), .B2(G150), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G303), .A2(new_n795), .B1(new_n775), .B2(G311), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT105), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT106), .B(G317), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n252), .B1(new_n792), .B2(new_n1035), .C1(new_n777), .C2(new_n411), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G97), .B2(new_n810), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n812), .A2(G116), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT46), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G283), .A2(new_n782), .B1(new_n797), .B2(G294), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1034), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1033), .A2(KEYINPUT105), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1032), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT47), .Z(new_n1044));
  OAI211_X1 g0844(.A(new_n768), .B(new_n1025), .C1(new_n1044), .C2(new_n859), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n978), .A2(new_n828), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1024), .A2(new_n1048), .ZN(G387));
  NAND2_X1  g0849(.A1(new_n1010), .A2(new_n767), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n202), .A2(new_n804), .B1(new_n803), .B2(new_n807), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n281), .B2(new_n797), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n787), .A2(new_n218), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n269), .B1(new_n792), .B2(new_n851), .C1(new_n477), .C2(new_n790), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n575), .C2(new_n778), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1052), .B(new_n1055), .C1(new_n258), .C2(new_n783), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G303), .A2(new_n782), .B1(new_n797), .B2(G311), .ZN(new_n1057));
  INV_X1    g0857(.A(G322), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n803), .C1(new_n804), .C2(new_n1035), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G294), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n777), .A2(new_n791), .B1(new_n787), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(KEYINPUT49), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n792), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n269), .B1(new_n1066), .B2(G326), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(new_n479), .C2(new_n790), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT49), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n771), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n714), .B(new_n290), .C1(new_n258), .C2(new_n218), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT107), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n399), .A2(G50), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT50), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n822), .B1(new_n231), .B2(new_n290), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(G107), .B2(new_n207), .C1(new_n714), .C2(new_n818), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n769), .B1(new_n1079), .B2(new_n829), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n828), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1071), .B(new_n1080), .C1(new_n706), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT104), .B1(new_n1010), .B2(new_n759), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1006), .B(new_n758), .C1(new_n1009), .C2(new_n1002), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n716), .B1(new_n1010), .B2(new_n759), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1050), .B(new_n1082), .C1(new_n1085), .C2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1021), .A2(new_n1019), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n717), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT110), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n1088), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1092), .B1(new_n1091), .B2(new_n1088), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1089), .A2(new_n767), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n243), .A2(new_n823), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n829), .B1(new_n477), .B2(new_n207), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n768), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT108), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G150), .A2(new_n775), .B1(new_n795), .B2(G159), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  OAI22_X1  g0903(.A1(new_n777), .A2(new_n218), .B1(new_n787), .B2(new_n258), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n252), .B1(new_n1066), .B2(G143), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n545), .B2(new_n790), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(G50), .C2(new_n797), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1107), .C1(new_n399), .C2(new_n783), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G311), .A2(new_n795), .B1(new_n775), .B2(G317), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n782), .A2(G294), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n777), .A2(new_n479), .B1(new_n787), .B2(new_n791), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n252), .B1(new_n792), .B2(new_n1058), .C1(new_n411), .C2(new_n790), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(new_n797), .C2(G303), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1101), .B1(new_n984), .B2(new_n1081), .C1(new_n1118), .C2(new_n859), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1097), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1096), .A2(new_n1121), .ZN(G390));
  AOI21_X1  g0922(.A(KEYINPUT111), .B1(new_n906), .B2(new_n933), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n904), .B1(new_n863), .B2(new_n899), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT111), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n933), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n924), .A2(new_n927), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n930), .A2(KEYINPUT39), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n924), .A2(new_n928), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n841), .A2(new_n418), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n730), .A2(new_n702), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n899), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1126), .B1(new_n1135), .B2(new_n905), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n842), .A2(G330), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n753), .B2(new_n755), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n905), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1131), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n931), .A2(new_n1128), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1138), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n944), .A2(new_n905), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n937), .A2(new_n648), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n448), .A2(new_n944), .A3(G330), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT112), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT112), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n960), .A2(new_n1149), .A3(G330), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1146), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n905), .B1(new_n756), .B2(new_n1143), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1138), .B(new_n904), .C1(new_n755), .C2(new_n943), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n900), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n904), .B1(new_n958), .B2(new_n1138), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1135), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1140), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT113), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1151), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n717), .B1(new_n1145), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1131), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1144), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1144), .B1(new_n905), .B2(new_n1139), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1135), .B1(new_n905), .B2(new_n1139), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n900), .A2(new_n1167), .B1(new_n1168), .B2(new_n1155), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1149), .B1(new_n960), .B2(G330), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1147), .A2(KEYINPUT112), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n938), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT113), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1151), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1166), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1163), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n931), .A2(new_n826), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n837), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n768), .B1(new_n281), .B2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n477), .A2(new_n783), .B1(new_n804), .B2(new_n479), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G107), .B2(new_n797), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n790), .A2(new_n258), .B1(new_n792), .B2(new_n1062), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT116), .Z(new_n1184));
  OAI221_X1 g0984(.A(new_n252), .B1(new_n787), .B2(new_n545), .C1(new_n777), .C2(new_n218), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n775), .B2(G283), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n782), .A2(new_n1189), .B1(G159), .B2(new_n778), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n850), .B2(new_n798), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT114), .ZN(new_n1192));
  INV_X1    g0992(.A(G125), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n269), .B1(new_n792), .B2(new_n1193), .C1(new_n202), .C2(new_n790), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT115), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT53), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n787), .B2(new_n851), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n812), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n795), .A2(G132), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G128), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1195), .B(new_n1199), .C1(new_n1200), .C2(new_n803), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1187), .B1(new_n1192), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT117), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n859), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1180), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1166), .A2(new_n767), .B1(new_n1178), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1177), .A2(new_n1207), .ZN(G378));
  INV_X1    g1008(.A(new_n392), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n686), .A2(new_n377), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  OR3_X1    g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n826), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n768), .B1(G50), .B2(new_n1179), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G50), .B1(new_n248), .B2(new_n289), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n269), .B2(G41), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n289), .B(new_n252), .C1(new_n792), .C2(new_n791), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n790), .A2(new_n257), .ZN(new_n1225));
  OR4_X1    g1025(.A1(new_n1026), .A2(new_n1224), .A3(new_n1053), .A4(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G97), .A2(new_n797), .B1(new_n795), .B2(G107), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n479), .B2(new_n803), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n575), .C2(new_n782), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1223), .B1(new_n1229), .B2(KEYINPUT58), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(KEYINPUT58), .B2(new_n1229), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G33), .B(G41), .C1(new_n1066), .C2(G124), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n795), .A2(G128), .B1(new_n812), .B2(new_n1189), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT118), .Z(new_n1234));
  OAI22_X1  g1034(.A1(new_n803), .A2(new_n1193), .B1(new_n851), .B2(new_n777), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n854), .A2(new_n798), .B1(new_n783), .B2(new_n850), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT59), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1232), .B1(new_n807), .B2(new_n790), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1231), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1221), .B1(new_n1241), .B2(new_n771), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n907), .B1(new_n1244), .B2(new_n1126), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n679), .B1(new_n952), .B2(new_n953), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n951), .A3(new_n1218), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n947), .B1(new_n928), .B2(new_n929), .ZN(new_n1248));
  OAI21_X1  g1048(.A(G330), .B1(new_n1248), .B2(KEYINPUT40), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT40), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n924), .B2(new_n928), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1219), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1245), .A2(new_n1247), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1244), .A2(new_n1126), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1252), .A2(new_n1247), .B1(new_n1254), .B2(new_n908), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1243), .B1(new_n1256), .B2(new_n766), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT57), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1172), .B1(new_n1166), .B2(new_n1175), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1256), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1218), .B1(new_n1246), .B2(new_n951), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1249), .A2(new_n1251), .A3(new_n1219), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n934), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1245), .A2(new_n1247), .A3(new_n1252), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1151), .B1(new_n1145), .B2(new_n1162), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n717), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1257), .B1(new_n1260), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(G375));
  NAND2_X1  g1069(.A1(new_n904), .A2(new_n826), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT119), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n252), .B1(new_n792), .B2(new_n451), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G77), .B2(new_n810), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n778), .A2(new_n575), .B1(new_n812), .B2(G97), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n783), .C2(new_n411), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(G116), .A2(new_n797), .B1(new_n795), .B2(G283), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1062), .B2(new_n803), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(G132), .A2(new_n775), .B1(new_n782), .B2(G150), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n798), .B2(new_n1188), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n777), .A2(new_n202), .B1(new_n787), .B2(new_n807), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n269), .B1(new_n792), .B2(new_n1200), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1280), .A2(new_n1225), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n804), .B2(new_n850), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1275), .A2(new_n1277), .B1(new_n1279), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT120), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n859), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1285), .B2(new_n1284), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n769), .B1(new_n258), .B2(new_n837), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1158), .A2(new_n767), .B1(new_n1271), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1291), .A2(new_n997), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1292), .B2(new_n1175), .ZN(G381));
  NOR2_X1   g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  INV_X1    g1094(.A(G378), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(G381), .A2(G384), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G387), .A2(G390), .A3(new_n1297), .A4(G375), .ZN(new_n1298));
  XOR2_X1   g1098(.A(new_n1298), .B(KEYINPUT121), .Z(G407));
  NAND3_X1  g1099(.A1(new_n1268), .A2(new_n687), .A3(new_n1295), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(G407), .A2(G213), .A3(new_n1300), .ZN(G409));
  XNOR2_X1  g1101(.A(G393), .B(new_n835), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n758), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n766), .B1(new_n1304), .B2(new_n997), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1047), .B1(new_n1305), .B2(new_n996), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G390), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT110), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1093), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1120), .B1(new_n1309), .B2(new_n1090), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(G387), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1303), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1306), .A2(G390), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1310), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1302), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1243), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1318), .A2(KEYINPUT123), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n766), .B1(new_n1318), .B2(KEYINPUT123), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OR3_X1    g1121(.A1(new_n1259), .A2(new_n1256), .A3(new_n997), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G378), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1317), .B1(new_n1318), .B2(new_n767), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n716), .B1(new_n1259), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT57), .B1(new_n1266), .B2(new_n1318), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G378), .B(new_n1325), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT122), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT122), .B1(new_n1268), .B2(G378), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1324), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(G213), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(G343), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1173), .A2(KEYINPUT60), .A3(new_n1174), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1291), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(KEYINPUT124), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1337), .A2(new_n1341), .A3(new_n1338), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n717), .B1(new_n1291), .B2(KEYINPUT60), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1340), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT125), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1343), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1346), .B1(new_n1339), .B2(KEYINPUT124), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT125), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(new_n1348), .A3(new_n1342), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1345), .A2(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(G384), .B1(new_n1350), .B2(new_n1290), .ZN(new_n1351));
  INV_X1    g1151(.A(G384), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1290), .ZN(new_n1353));
  AOI211_X1 g1153(.A(new_n1352), .B(new_n1353), .C1(new_n1345), .C2(new_n1349), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1351), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1333), .A2(new_n1336), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(KEYINPUT126), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT126), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1333), .A2(new_n1355), .A3(new_n1358), .A4(new_n1336), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT62), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1360));
  AND4_X1   g1160(.A1(new_n1348), .A2(new_n1340), .A3(new_n1342), .A4(new_n1343), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1348), .B1(new_n1347), .B2(new_n1342), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1290), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n1352), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1350), .A2(G384), .A3(new_n1290), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1335), .A2(G2897), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  AND3_X1   g1167(.A1(new_n1364), .A2(new_n1365), .A3(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1367), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1268), .A2(KEYINPUT122), .A3(G378), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1323), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  OAI22_X1  g1172(.A1(new_n1368), .A2(new_n1369), .B1(new_n1372), .B2(new_n1335), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT61), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT62), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1376));
  NOR3_X1   g1176(.A1(new_n1372), .A2(new_n1376), .A3(new_n1335), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1373), .B(new_n1374), .C1(new_n1375), .C2(new_n1377), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1316), .B1(new_n1360), .B2(new_n1378), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1312), .A2(new_n1374), .A3(new_n1315), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1380), .B1(KEYINPUT63), .B2(new_n1377), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1355), .A2(new_n1367), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT127), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1376), .A2(new_n1366), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1382), .A2(new_n1383), .A3(new_n1384), .ZN(new_n1385));
  OAI21_X1  g1185(.A(KEYINPUT127), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1386));
  OAI211_X1 g1186(.A(new_n1385), .B(new_n1386), .C1(new_n1335), .C2(new_n1372), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT63), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1357), .A2(new_n1388), .A3(new_n1359), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1381), .A2(new_n1387), .A3(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1379), .A2(new_n1390), .ZN(G405));
  AOI22_X1  g1191(.A1(new_n1370), .A2(new_n1371), .B1(new_n1295), .B2(G375), .ZN(new_n1392));
  XNOR2_X1  g1192(.A(new_n1392), .B(new_n1376), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(new_n1393), .B(new_n1316), .ZN(G402));
endmodule


