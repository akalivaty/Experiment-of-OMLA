

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U328 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U329 ( .A(n453), .B(n452), .ZN(n567) );
  AND2_X1 U330 ( .A1(n472), .A2(n550), .ZN(n296) );
  XOR2_X1 U331 ( .A(G85GAT), .B(KEYINPUT70), .Z(n297) );
  XOR2_X1 U332 ( .A(n322), .B(n362), .Z(n298) );
  INV_X1 U333 ( .A(KEYINPUT110), .ZN(n385) );
  XNOR2_X1 U334 ( .A(n386), .B(n385), .ZN(n387) );
  INV_X1 U335 ( .A(KEYINPUT73), .ZN(n326) );
  XNOR2_X1 U336 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U337 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U338 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U339 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n384) );
  XNOR2_X1 U340 ( .A(n579), .B(n384), .ZN(n506) );
  XOR2_X1 U341 ( .A(n334), .B(n333), .Z(n584) );
  NOR2_X1 U342 ( .A1(n467), .A2(n456), .ZN(n564) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U344 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(G71GAT), .B(KEYINPUT81), .Z(n300) );
  XNOR2_X1 U346 ( .A(KEYINPUT80), .B(KEYINPUT20), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n310) );
  XOR2_X1 U348 ( .A(KEYINPUT0), .B(KEYINPUT75), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT76), .B(G120GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(G113GAT), .B(n303), .Z(n437) );
  XOR2_X1 U352 ( .A(KEYINPUT77), .B(G99GAT), .Z(n305) );
  XOR2_X1 U353 ( .A(G43GAT), .B(G134GAT), .Z(n345) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .Z(n322) );
  XNOR2_X1 U355 ( .A(n345), .B(n322), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U357 ( .A(n437), .B(n306), .Z(n308) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n318) );
  XOR2_X1 U361 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n312) );
  XNOR2_X1 U362 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U364 ( .A(n313), .B(KEYINPUT19), .Z(n315) );
  XNOR2_X1 U365 ( .A(G190GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U367 ( .A(G169GAT), .B(G176GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n409) );
  XOR2_X2 U369 ( .A(n318), .B(n409), .Z(n532) );
  INV_X1 U370 ( .A(n532), .ZN(n467) );
  XNOR2_X1 U371 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n414) );
  XOR2_X1 U372 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n320) );
  XNOR2_X1 U373 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n334) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(G1GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n321), .B(KEYINPUT67), .ZN(n362) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n298), .B(n323), .ZN(n329) );
  XOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .Z(n325) );
  XNOR2_X1 U380 ( .A(G71GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n372) );
  XNOR2_X1 U382 ( .A(n372), .B(KEYINPUT15), .ZN(n327) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G155GAT), .Z(n419) );
  XOR2_X1 U384 ( .A(n330), .B(n419), .Z(n332) );
  XNOR2_X1 U385 ( .A(G183GAT), .B(G211GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n336) );
  XNOR2_X1 U388 ( .A(G92GAT), .B(KEYINPUT72), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n349) );
  XNOR2_X1 U390 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n337), .B(KEYINPUT7), .ZN(n358) );
  XOR2_X1 U392 ( .A(n358), .B(KEYINPUT11), .Z(n339) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G106GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n297), .B(n340), .ZN(n373) );
  XOR2_X1 U397 ( .A(n341), .B(n373), .Z(n343) );
  XOR2_X1 U398 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U399 ( .A(G36GAT), .B(G218GAT), .Z(n404) );
  XNOR2_X1 U400 ( .A(n423), .B(n404), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U402 ( .A(n344), .B(KEYINPUT9), .Z(n347) );
  XNOR2_X1 U403 ( .A(G190GAT), .B(n345), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n390) );
  INV_X1 U406 ( .A(n390), .ZN(n560) );
  XOR2_X1 U407 ( .A(KEYINPUT36), .B(KEYINPUT98), .Z(n350) );
  XNOR2_X1 U408 ( .A(n560), .B(n350), .ZN(n588) );
  NOR2_X1 U409 ( .A1(n584), .A2(n588), .ZN(n351) );
  XNOR2_X1 U410 ( .A(KEYINPUT45), .B(n351), .ZN(n383) );
  XOR2_X1 U411 ( .A(G22GAT), .B(G141GAT), .Z(n353) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G113GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U414 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n355) );
  XNOR2_X1 U415 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n368) );
  XOR2_X1 U418 ( .A(n358), .B(KEYINPUT29), .Z(n360) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(G169GAT), .B(n361), .ZN(n366) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G36GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(G43GAT), .B(n362), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n551) );
  XOR2_X1 U427 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n370) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U430 ( .A(n371), .B(KEYINPUT71), .Z(n375) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U433 ( .A(KEYINPUT69), .B(KEYINPUT33), .Z(n377) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G120GAT), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U436 ( .A(n379), .B(n378), .Z(n381) );
  XOR2_X1 U437 ( .A(G204GAT), .B(G148GAT), .Z(n426) );
  XOR2_X1 U438 ( .A(G92GAT), .B(G64GAT), .Z(n397) );
  XNOR2_X1 U439 ( .A(n426), .B(n397), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n579) );
  NOR2_X1 U441 ( .A1(n551), .A2(n579), .ZN(n382) );
  NAND2_X1 U442 ( .A1(n383), .A2(n382), .ZN(n395) );
  XNOR2_X1 U443 ( .A(n584), .B(KEYINPUT109), .ZN(n565) );
  INV_X1 U444 ( .A(n551), .ZN(n571) );
  NOR2_X1 U445 ( .A1(n571), .A2(n506), .ZN(n388) );
  XNOR2_X1 U446 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n386) );
  NOR2_X1 U447 ( .A1(n565), .A2(n389), .ZN(n391) );
  NAND2_X1 U448 ( .A1(n391), .A2(n390), .ZN(n393) );
  XOR2_X1 U449 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n392) );
  NAND2_X1 U450 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT48), .B(n396), .ZN(n548) );
  XOR2_X1 U452 ( .A(KEYINPUT92), .B(n397), .Z(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n399) );
  XNOR2_X1 U454 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(n400), .ZN(n433) );
  INV_X1 U457 ( .A(n433), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n401), .B(G204GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT91), .B(n404), .Z(n406) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n412) );
  INV_X1 U464 ( .A(n409), .ZN(n410) );
  XNOR2_X1 U465 ( .A(G8GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n522) );
  AND2_X1 U467 ( .A1(n548), .A2(n522), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n568) );
  INV_X1 U469 ( .A(n568), .ZN(n454) );
  XOR2_X1 U470 ( .A(KEYINPUT87), .B(KEYINPUT83), .Z(n416) );
  XNOR2_X1 U471 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n431) );
  XOR2_X1 U473 ( .A(KEYINPUT24), .B(G78GAT), .Z(n418) );
  XNOR2_X1 U474 ( .A(G218GAT), .B(G106GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n429) );
  XOR2_X1 U477 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n422) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n436) );
  XOR2_X1 U480 ( .A(n436), .B(n423), .Z(n425) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n431), .B(n430), .Z(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n472) );
  XOR2_X1 U487 ( .A(KEYINPUT89), .B(G57GAT), .Z(n435) );
  XNOR2_X1 U488 ( .A(G1GAT), .B(G155GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n439) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n453) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n447) );
  XOR2_X1 U495 ( .A(G85GAT), .B(G148GAT), .Z(n443) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(G127GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U498 ( .A(G134GAT), .B(G162GAT), .Z(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n449) );
  XNOR2_X1 U502 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U505 ( .A(n567), .ZN(n550) );
  NAND2_X1 U506 ( .A1(n454), .A2(n296), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT55), .B(n455), .Z(n456) );
  NAND2_X1 U508 ( .A1(n564), .A2(n560), .ZN(n458) );
  NAND2_X1 U509 ( .A1(n564), .A2(n551), .ZN(n460) );
  XNOR2_X1 U510 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n460), .B(n459), .ZN(G1348GAT) );
  INV_X1 U512 ( .A(n506), .ZN(n553) );
  NAND2_X1 U513 ( .A1(n564), .A2(n553), .ZN(n464) );
  XOR2_X1 U514 ( .A(G176GAT), .B(KEYINPUT121), .Z(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  NOR2_X1 U518 ( .A1(n579), .A2(n571), .ZN(n494) );
  XNOR2_X1 U519 ( .A(n522), .B(KEYINPUT93), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT27), .ZN(n470) );
  XOR2_X1 U521 ( .A(n472), .B(KEYINPUT28), .Z(n527) );
  NOR2_X1 U522 ( .A1(n470), .A2(n527), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n567), .A2(n466), .ZN(n534) );
  XOR2_X1 U524 ( .A(KEYINPUT82), .B(n467), .Z(n468) );
  NOR2_X1 U525 ( .A1(n534), .A2(n468), .ZN(n479) );
  NOR2_X1 U526 ( .A1(n532), .A2(n472), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT26), .B(n469), .Z(n569) );
  NOR2_X1 U528 ( .A1(n470), .A2(n569), .ZN(n547) );
  NAND2_X1 U529 ( .A1(n532), .A2(n522), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT94), .B(n471), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U532 ( .A(n474), .B(KEYINPUT25), .Z(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT95), .B(n475), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n547), .A2(n476), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n567), .A2(n477), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n491) );
  NOR2_X1 U537 ( .A1(n560), .A2(n584), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U539 ( .A1(n491), .A2(n481), .ZN(n507) );
  AND2_X1 U540 ( .A1(n494), .A2(n507), .ZN(n489) );
  NAND2_X1 U541 ( .A1(n489), .A2(n567), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n489), .A2(n522), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U547 ( .A1(n489), .A2(n532), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n488) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT96), .Z(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n489), .A2(n527), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n498) );
  NOR2_X1 U554 ( .A1(n491), .A2(n588), .ZN(n492) );
  NAND2_X1 U555 ( .A1(n584), .A2(n492), .ZN(n493) );
  XNOR2_X1 U556 ( .A(KEYINPUT37), .B(n493), .ZN(n518) );
  NAND2_X1 U557 ( .A1(n518), .A2(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT38), .B(KEYINPUT99), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n567), .A2(n503), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n503), .A2(n522), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n532), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(KEYINPUT40), .ZN(n502) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  XOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT101), .Z(n505) );
  NAND2_X1 U569 ( .A1(n527), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  NOR2_X1 U571 ( .A1(n551), .A2(n506), .ZN(n519) );
  AND2_X1 U572 ( .A1(n519), .A2(n507), .ZN(n514) );
  NAND2_X1 U573 ( .A1(n514), .A2(n567), .ZN(n511) );
  XOR2_X1 U574 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n514), .A2(n522), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n532), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U583 ( .A1(n514), .A2(n527), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT105), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n567), .A2(n528), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n522), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT106), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  XOR2_X1 U593 ( .A(G99GAT), .B(KEYINPUT107), .Z(n526) );
  NAND2_X1 U594 ( .A1(n528), .A2(n532), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n530) );
  NAND2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n531), .Z(G1339GAT) );
  NAND2_X1 U600 ( .A1(n532), .A2(n548), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n542), .A2(n551), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U605 ( .A1(n542), .A2(n553), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U609 ( .A1(n542), .A2(n565), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U613 ( .A1(n542), .A2(n560), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT115), .Z(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n551), .A2(n561), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n555) );
  NAND2_X1 U622 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  INV_X1 U626 ( .A(n584), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT118), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  OR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n580) );
  INV_X1 U636 ( .A(n580), .ZN(n587) );
  NOR2_X1 U637 ( .A1(n587), .A2(n571), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT122), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(n574), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

