//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(KEYINPUT3), .A3(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n463), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n470), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n463), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n476), .A2(G2105), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(KEYINPUT68), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI221_X1 g060(.A(new_n478), .B1(new_n479), .B2(new_n480), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n463), .A2(G138), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n461), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n469), .A2(new_n470), .A3(new_n490), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n493), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n470), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT6), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(KEYINPUT72), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n504), .B(KEYINPUT6), .C1(new_n505), .C2(KEYINPUT72), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n508), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n516), .A2(G62), .ZN(new_n519));
  AND2_X1   g094(.A1(G75), .A2(G543), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n513), .A2(new_n518), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(G76), .A2(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n505), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  INV_X1    g102(.A(new_n517), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(G89), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n526), .B1(new_n511), .B2(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n516), .B(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G63), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n524), .A2(new_n525), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n505), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(new_n531), .A2(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n505), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n511), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AND2_X1   g117(.A1(new_n531), .A2(G56), .ZN(new_n543));
  AND2_X1   g118(.A1(G68), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n512), .A2(G43), .B1(G81), .B2(new_n517), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n511), .B2(new_n554), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n517), .A2(G91), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(G65), .Z(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(new_n516), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n505), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  NAND2_X1  g139(.A1(new_n512), .A2(G49), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n517), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT77), .Z(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n514), .B2(new_n515), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n508), .A2(G48), .A3(G543), .A4(new_n509), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n508), .A2(G86), .A3(new_n509), .A4(new_n516), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n512), .A2(G47), .B1(G85), .B2(new_n517), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n505), .B2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n516), .A2(G66), .ZN(new_n581));
  AND2_X1   g156(.A1(G79), .A2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G54), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT10), .B1(new_n517), .B2(G92), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n583), .B1(new_n584), .B2(new_n511), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n580), .B1(G868), .B2(new_n589), .ZN(G284));
  OAI21_X1  g165(.A(new_n580), .B1(G868), .B2(new_n589), .ZN(G321));
  NAND2_X1  g166(.A1(G286), .A2(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n557), .A2(new_n561), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(G868), .ZN(G297));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(G868), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g176(.A(new_n484), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G135), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n477), .A2(G123), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT78), .Z(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  INV_X1    g182(.A(G111), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n606), .A2(new_n607), .B1(new_n608), .B2(G2105), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n607), .B2(new_n606), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n603), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(G2096), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n472), .A2(new_n461), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(G156));
  XOR2_X1   g193(.A(G2451), .B(G2454), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT16), .ZN(new_n620));
  XNOR2_X1  g195(.A(G1341), .B(G1348), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(new_n625), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n622), .B(new_n628), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(G14), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n630), .ZN(G401));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n635), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n636), .A2(new_n637), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2096), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1956), .B(G2474), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n650), .A2(new_n652), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n655), .A3(new_n653), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n658), .B(new_n661), .C1(new_n655), .C2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  MUX2_X1   g243(.A(G6), .B(G305), .S(G16), .Z(new_n669));
  XOR2_X1   g244(.A(KEYINPUT32), .B(G1981), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n672), .A2(KEYINPUT85), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(KEYINPUT85), .ZN(new_n674));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G23), .ZN(new_n676));
  INV_X1    g251(.A(G288), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT33), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(G22), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G166), .B2(new_n675), .ZN(new_n683));
  INV_X1    g258(.A(G1971), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND4_X1  g260(.A1(new_n673), .A2(new_n674), .A3(new_n681), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT87), .Z(new_n687));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n477), .A2(G119), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n463), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n602), .B2(G131), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT84), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G29), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G25), .B2(G29), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  MUX2_X1   g276(.A(G24), .B(G290), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n689), .A2(new_n690), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT36), .Z(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G35), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G162), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G2090), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT91), .B1(G16), .B2(G21), .ZN(new_n713));
  NAND2_X1  g288(.A1(G168), .A2(G16), .ZN(new_n714));
  MUX2_X1   g289(.A(KEYINPUT91), .B(new_n713), .S(new_n714), .Z(new_n715));
  INV_X1    g290(.A(G1966), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n707), .A2(G32), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT26), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n477), .A2(G129), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n720), .B(new_n721), .C1(G105), .C2(new_n472), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n602), .A2(G141), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n707), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT27), .B(G1996), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G171), .A2(new_n675), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G5), .B2(new_n675), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n707), .B2(new_n611), .ZN(new_n733));
  AND2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n707), .B1(KEYINPUT24), .B2(G34), .ZN(new_n735));
  OAI22_X1  g310(.A1(G160), .A2(new_n707), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n730), .A2(new_n731), .B1(G2084), .B2(new_n736), .ZN(new_n737));
  NOR4_X1   g312(.A1(new_n717), .A2(new_n728), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n675), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT23), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n593), .B2(new_n675), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n707), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n707), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G2078), .Z(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G19), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n548), .B2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1341), .Z(new_n749));
  XOR2_X1   g324(.A(KEYINPUT31), .B(G11), .Z(new_n750));
  AND2_X1   g325(.A1(new_n736), .A2(G2084), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT92), .B(G28), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT30), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(KEYINPUT30), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n750), .B(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT25), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(new_n463), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n758), .B1(new_n760), .B2(KEYINPUT90), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n761), .B1(KEYINPUT90), .B2(new_n760), .C1(new_n484), .C2(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G33), .B(new_n763), .S(G29), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n707), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n602), .A2(G140), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n463), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n477), .A2(G128), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT89), .B(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n589), .B2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT88), .B(G1348), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n756), .A2(new_n765), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n738), .A2(new_n743), .A3(new_n746), .A4(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n706), .A2(new_n712), .A3(new_n782), .ZN(G311));
  INV_X1    g358(.A(G311), .ZN(G150));
  NAND2_X1  g359(.A1(new_n531), .A2(G67), .ZN(new_n785));
  NAND2_X1  g360(.A1(G80), .A2(G543), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G651), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n512), .A2(G55), .B1(G93), .B2(new_n517), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n547), .B1(new_n790), .B2(KEYINPUT94), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(KEYINPUT94), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n589), .A2(G559), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n795), .B(new_n796), .Z(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT39), .ZN(new_n798));
  INV_X1    g373(.A(G860), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(KEYINPUT39), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n790), .A2(new_n799), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT37), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(G145));
  NAND2_X1  g379(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n724), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n477), .A2(G130), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n463), .A2(G118), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n602), .B2(G142), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n615), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n806), .B(new_n812), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n493), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n814));
  AOI21_X1  g389(.A(KEYINPUT70), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n491), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n499), .A2(KEYINPUT96), .A3(new_n501), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT96), .B1(new_n499), .B2(new_n501), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n773), .B(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n696), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n813), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n611), .B(G160), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n487), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  AOI21_X1  g402(.A(G37), .B1(new_n823), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g405(.A(new_n793), .B(new_n598), .ZN(new_n831));
  NAND2_X1  g406(.A1(G299), .A2(new_n589), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n588), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT99), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT41), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT100), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n834), .B(KEYINPUT41), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(KEYINPUT100), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n836), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT42), .ZN(new_n842));
  XOR2_X1   g417(.A(G288), .B(KEYINPUT101), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G305), .ZN(new_n844));
  XNOR2_X1  g419(.A(G290), .B(G303), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n842), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G868), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G868), .B2(new_n790), .ZN(G295));
  OAI21_X1  g424(.A(new_n848), .B1(G868), .B2(new_n790), .ZN(G331));
  XNOR2_X1  g425(.A(G168), .B(G171), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n793), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT102), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT102), .ZN(new_n855));
  INV_X1    g430(.A(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n834), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n846), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n854), .A2(new_n846), .A3(new_n855), .A4(new_n857), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT43), .ZN(new_n864));
  INV_X1    g439(.A(new_n862), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT43), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n846), .B1(new_n856), .B2(new_n835), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n852), .A2(new_n839), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(KEYINPUT44), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n862), .A2(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT103), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n862), .A2(new_n876), .A3(new_n869), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(KEYINPUT43), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n866), .A2(new_n861), .A3(new_n860), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n872), .A2(new_n880), .ZN(G397));
  INV_X1    g456(.A(G1384), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n502), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n499), .A2(KEYINPUT96), .A3(new_n501), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n882), .B1(new_n498), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(G160), .A2(G40), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G1996), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n724), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G2067), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n773), .B(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n894), .A2(new_n696), .A3(new_n896), .A4(new_n699), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n768), .A2(new_n895), .A3(new_n772), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n696), .B(new_n699), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n896), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(KEYINPUT126), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n892), .A2(G1986), .A3(G290), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT48), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(KEYINPUT126), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n891), .A2(new_n893), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT46), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n896), .A2(new_n725), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n892), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT125), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n908), .B1(KEYINPUT47), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(KEYINPUT47), .B2(new_n913), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT63), .ZN(new_n916));
  AND2_X1   g491(.A1(G160), .A2(G40), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n820), .A2(new_n917), .A3(new_n882), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n565), .A2(G1976), .A3(new_n566), .A4(new_n567), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(G8), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT52), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n920), .B2(KEYINPUT52), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G305), .A2(G1981), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(G1981), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n573), .A2(new_n574), .A3(new_n575), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(G305), .A2(KEYINPUT106), .A3(G1981), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT49), .ZN(new_n932));
  INV_X1    g507(.A(G8), .ZN(new_n933));
  AOI21_X1  g508(.A(G1384), .B1(new_n816), .B2(new_n819), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n917), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT49), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n936), .A3(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n677), .B2(G1976), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n920), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n924), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G2090), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT50), .B1(new_n820), .B2(new_n882), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  INV_X1    g520(.A(new_n502), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n945), .B(G1384), .C1(new_n816), .C2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n943), .B(new_n917), .C1(new_n944), .C2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n888), .A2(G1384), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n498), .B2(new_n886), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n816), .B2(new_n946), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n917), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n684), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n933), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT104), .B(KEYINPUT55), .ZN(new_n955));
  AND3_X1   g530(.A1(G303), .A2(G8), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(G303), .B2(G8), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n917), .B1(new_n934), .B2(new_n945), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n951), .A2(new_n945), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT107), .B(new_n917), .C1(new_n934), .C2(new_n945), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n943), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n933), .B1(new_n966), .B2(new_n953), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n942), .B(new_n960), .C1(new_n967), .C2(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n816), .A2(new_n946), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n890), .B1(new_n969), .B2(new_n949), .ZN(new_n970));
  AOI21_X1  g545(.A(G1966), .B1(new_n889), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n890), .A2(G2084), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n887), .A2(new_n945), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n951), .A2(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n977), .A2(new_n933), .A3(G286), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n916), .B1(new_n968), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n954), .A2(new_n959), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n940), .A2(new_n920), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(new_n938), .C1(new_n922), .C2(new_n923), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n954), .A2(new_n959), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(KEYINPUT63), .A3(new_n978), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n938), .A2(new_n988), .A3(new_n677), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n928), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n942), .A2(new_n981), .B1(new_n990), .B2(new_n935), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT62), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT116), .B1(new_n971), .B2(new_n976), .ZN(new_n994));
  INV_X1    g569(.A(new_n949), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n917), .B1(G164), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n820), .B2(new_n882), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n716), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n972), .B1(new_n944), .B2(new_n947), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n933), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G168), .A2(new_n933), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT117), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT51), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1003), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1006), .B(new_n1007), .C1(new_n977), .C2(new_n933), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n994), .B2(new_n1001), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n993), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n966), .A2(new_n953), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n958), .B1(new_n1013), .B2(new_n933), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n917), .B1(new_n944), .B2(new_n947), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT118), .B(G1961), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(G2078), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n889), .A2(new_n970), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n952), .B2(G2078), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G171), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n984), .A2(new_n1014), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1010), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n993), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1012), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g604(.A(KEYINPUT62), .B(new_n1010), .C1(new_n1005), .C2(new_n1008), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT123), .B1(new_n1030), .B2(new_n1025), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n992), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT122), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n971), .A2(new_n976), .A3(KEYINPUT116), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n999), .B1(new_n998), .B2(new_n1000), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1004), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1006), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1008), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1011), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n968), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n471), .A2(KEYINPUT119), .A3(new_n473), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1019), .A2(G40), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n464), .B(new_n1045), .C1(new_n474), .C2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n889), .A2(new_n950), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1017), .A2(new_n1021), .A3(G301), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1023), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT120), .B(KEYINPUT54), .C1(new_n1023), .C2(new_n1049), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1017), .A2(new_n1021), .A3(new_n1048), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1054), .B2(G171), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1017), .A2(new_n1021), .A3(G301), .A4(new_n1020), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1052), .A2(new_n1053), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1033), .B1(new_n1042), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1026), .A2(new_n968), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT54), .B1(new_n1023), .B2(new_n1049), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(new_n1043), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1054), .A2(G171), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(KEYINPUT54), .A3(new_n1057), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT121), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1062), .A2(new_n1064), .A3(KEYINPUT122), .A4(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT56), .B(G2072), .Z(new_n1069));
  NOR2_X1   g644(.A1(new_n952), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n742), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1073), .A3(new_n742), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n557), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n555), .A2(new_n1080), .A3(new_n556), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n561), .A2(KEYINPUT111), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n561), .A2(KEYINPUT111), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1079), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT112), .B(new_n1079), .C1(new_n1081), .C2(new_n1085), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1088), .B(new_n1089), .C1(new_n1079), .C2(G299), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n890), .B1(new_n974), .B2(new_n975), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1091), .A2(G1348), .B1(G2067), .B2(new_n918), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1078), .A2(new_n1090), .B1(new_n588), .B2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1070), .B(KEYINPUT113), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1077), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1090), .B(new_n1095), .C1(new_n1096), .C2(new_n1075), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1092), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n589), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1099), .B(new_n588), .C1(new_n1092), .C2(new_n1100), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1105), .A2(new_n1106), .B1(new_n1097), .B2(KEYINPUT61), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1097), .A2(KEYINPUT61), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n918), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n952), .B2(G1996), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT114), .A3(new_n548), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT59), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1098), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1061), .A2(new_n1068), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1032), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n900), .A2(new_n901), .ZN(new_n1118));
  XOR2_X1   g693(.A(G290), .B(G1986), .Z(new_n1119));
  AOI21_X1  g694(.A(new_n892), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT124), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1123), .B(new_n1120), .C1(new_n1032), .C2(new_n1116), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n915), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT127), .B(new_n915), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g704(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n871), .A2(new_n829), .A3(new_n1131), .ZN(G225));
  INV_X1    g706(.A(G225), .ZN(G308));
endmodule


