//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT67), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT67), .B1(new_n191), .B2(new_n193), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n195), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n197), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT11), .B1(new_n203), .B2(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n209), .B2(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n208), .A4(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n206), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .ZN(new_n227));
  OR2_X1    g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n234), .B(KEYINPUT1), .C1(new_n223), .C2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n234), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n225), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n239), .A3(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n210), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n209), .A2(G137), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n217), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n233), .A2(KEYINPUT30), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n231), .B1(new_n217), .B2(new_n219), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n217), .A2(new_n241), .A3(KEYINPUT66), .A4(new_n244), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n202), .B(new_n246), .C1(new_n251), .C2(KEYINPUT30), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT26), .B(G101), .Z(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G953), .ZN(new_n259));
  OR2_X1    g073(.A1(KEYINPUT68), .A2(G237), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT68), .A2(G237), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n257), .A2(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n255), .B(new_n263), .Z(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n202), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n233), .A2(new_n266), .A3(new_n245), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n252), .A2(KEYINPUT31), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT31), .B1(new_n252), .B2(new_n268), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n251), .B2(new_n266), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  INV_X1    g088(.A(new_n245), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n247), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n233), .A2(KEYINPUT71), .A3(new_n245), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n265), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n271), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n252), .A2(new_n268), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n252), .A2(KEYINPUT31), .A3(new_n268), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(new_n280), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n264), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n283), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n189), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT72), .B1(new_n271), .B2(new_n281), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n288), .A2(new_n283), .A3(new_n290), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n188), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT32), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n278), .A2(new_n299), .A3(new_n279), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n278), .B2(new_n279), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n202), .B1(new_n275), .B2(new_n247), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n279), .B1(new_n302), .B2(new_n267), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n252), .A2(new_n267), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT29), .B1(new_n307), .B2(new_n264), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n289), .B2(new_n264), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT75), .B(G902), .Z(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n294), .A2(new_n298), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G478), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(KEYINPUT15), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT97), .ZN(new_n317));
  INV_X1    g131(.A(G122), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G116), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n192), .A2(G122), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT94), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G107), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n192), .A2(G122), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(G116), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT94), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n223), .A2(G128), .ZN(new_n328));
  INV_X1    g142(.A(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G143), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G134), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n330), .A3(new_n209), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n319), .A2(KEYINPUT14), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n323), .A2(new_n324), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n335), .B(G107), .C1(new_n336), .C2(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n327), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT96), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT96), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n327), .A2(new_n334), .A3(new_n337), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n326), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n325), .B1(new_n323), .B2(new_n324), .ZN(new_n344));
  OAI21_X1  g158(.A(G107), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n327), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT13), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT13), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n223), .A3(G128), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n349), .A3(G134), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n346), .A2(new_n352), .A3(new_n333), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n342), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT9), .B(G234), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n357), .A2(new_n358), .A3(G953), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n342), .A2(new_n354), .A3(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n317), .B1(new_n363), .B2(new_n311), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n342), .A2(new_n354), .A3(new_n359), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n359), .B1(new_n342), .B2(new_n354), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n317), .B(new_n311), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n316), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT98), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n311), .B1(new_n365), .B2(new_n366), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n316), .B1(new_n371), .B2(KEYINPUT97), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n316), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(KEYINPUT97), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT98), .B1(new_n377), .B2(new_n372), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT92), .B(G143), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n262), .B2(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n260), .A2(new_n261), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n257), .A2(new_n259), .ZN(new_n383));
  NOR2_X1   g197(.A1(KEYINPUT92), .A2(G143), .ZN(new_n384));
  AND4_X1   g198(.A1(G214), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n208), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT17), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n383), .A3(G214), .ZN(new_n388));
  INV_X1    g202(.A(new_n380), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n262), .A2(G214), .A3(new_n384), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT17), .A4(G131), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G125), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT77), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G125), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n399), .A3(G140), .ZN(new_n400));
  INV_X1    g214(.A(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(KEYINPUT78), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT77), .B(G125), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n401), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT79), .A4(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n405), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n412), .A2(KEYINPUT16), .A3(G140), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n221), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(G146), .A3(new_n414), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n395), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G113), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(G104), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n390), .A2(new_n391), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n208), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n422), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT93), .A4(new_n425), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n403), .A2(new_n406), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G146), .ZN(new_n432));
  XOR2_X1   g246(.A(G125), .B(G140), .Z(new_n433));
  OR2_X1    g247(.A1(new_n433), .A2(G146), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n418), .A2(new_n421), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n386), .A2(new_n392), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n431), .B2(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n221), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n417), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n436), .ZN(new_n444));
  INV_X1    g258(.A(new_n421), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G475), .ZN(new_n448));
  INV_X1    g262(.A(G902), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G146), .B1(new_n411), .B2(new_n414), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n393), .A2(new_n394), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n221), .B(new_n413), .C1(new_n409), .C2(new_n410), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n436), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n456), .A2(new_n457), .A3(new_n445), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n421), .B1(new_n418), .B2(new_n436), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G475), .ZN(new_n461));
  NAND2_X1  g275(.A1(G234), .A2(G237), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n462), .A2(G952), .A3(new_n256), .ZN(new_n463));
  INV_X1    g277(.A(new_n383), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n310), .A3(new_n462), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT99), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G475), .B1(new_n437), .B2(new_n446), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n449), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n452), .A2(new_n461), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n379), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n231), .A2(new_n405), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n238), .A2(new_n240), .A3(new_n412), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n256), .A2(G224), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(new_n420), .B2(G107), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT82), .B(KEYINPUT3), .C1(new_n420), .C2(G107), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n420), .A2(KEYINPUT3), .A3(G107), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n420), .A2(G107), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G101), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n420), .A2(KEYINPUT3), .A3(G107), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n480), .B2(new_n479), .ZN(new_n488));
  INV_X1    g302(.A(G101), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n484), .A4(new_n482), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n490), .A3(KEYINPUT4), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n492), .A3(G101), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n493), .A3(new_n202), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G122), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n496), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n420), .B2(G107), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n322), .A2(KEYINPUT83), .A3(G104), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n484), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G101), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n485), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n489), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT67), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n194), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G116), .B(G119), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT67), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g326(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n196), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n494), .A2(new_n499), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n499), .B(KEYINPUT87), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n494), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT6), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n494), .A2(new_n516), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n518), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n478), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n497), .A2(new_n526), .A3(new_n498), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n497), .B2(new_n498), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT8), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT89), .B1(new_n507), .B2(new_n515), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n490), .A2(new_n504), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n513), .B1(new_n200), .B2(KEYINPUT5), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n196), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n513), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n540));
  OR3_X1    g354(.A1(new_n535), .A2(new_n196), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n533), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n494), .A2(new_n499), .A3(new_n516), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n477), .A2(KEYINPUT7), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n474), .B(new_n475), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n474), .B2(new_n544), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n548), .A2(new_n476), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n542), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G210), .B1(G237), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR4_X1   g366(.A1(new_n524), .A2(new_n550), .A3(G902), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n551), .B(KEYINPUT91), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n520), .A2(new_n523), .ZN(new_n556));
  INV_X1    g370(.A(new_n478), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n550), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n553), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n473), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT23), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n190), .B2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n329), .A2(KEYINPUT23), .A3(G119), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n571), .B(new_n572), .C1(G119), .C2(new_n329), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n568), .A2(KEYINPUT76), .B1(new_n573), .B2(G110), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n569), .B(new_n574), .C1(new_n453), .C2(new_n455), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n573), .A2(G110), .B1(new_n567), .B2(new_n566), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n417), .A2(new_n576), .A3(new_n434), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n383), .A2(G221), .A3(G234), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(new_n577), .A3(new_n581), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n311), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT25), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n358), .B1(new_n311), .B2(G234), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n583), .A2(new_n588), .A3(new_n311), .A4(new_n584), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n583), .A2(new_n584), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n587), .A2(G902), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n314), .A2(new_n565), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G469), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n217), .A2(new_n219), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT84), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n240), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n226), .A2(KEYINPUT84), .A3(new_n239), .A4(G128), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n239), .B1(G143), .B2(new_n221), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n225), .B1(new_n602), .B2(new_n329), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n507), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n535), .A2(new_n240), .A3(new_n238), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n507), .A2(KEYINPUT10), .A3(new_n241), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n491), .A2(new_n232), .A3(new_n493), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n598), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n383), .A2(G227), .ZN(new_n615));
  XNOR2_X1  g429(.A(G110), .B(G140), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n220), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(new_n614), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n597), .B(new_n311), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT85), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n614), .A2(KEYINPUT85), .A3(new_n617), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n617), .ZN(new_n628));
  INV_X1    g442(.A(new_n614), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n628), .B1(new_n609), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(new_n630), .A3(G469), .ZN(new_n631));
  NAND2_X1  g445(.A1(G469), .A2(G902), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n623), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(G221), .B1(new_n357), .B2(G902), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT81), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n596), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT100), .B(G101), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G3));
  AOI21_X1  g453(.A(new_n310), .B1(new_n295), .B2(new_n296), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n292), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n633), .A2(new_n635), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n595), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n452), .A2(new_n461), .A3(new_n471), .ZN(new_n646));
  INV_X1    g460(.A(new_n363), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT33), .B1(new_n647), .B2(KEYINPUT102), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n363), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n310), .A2(new_n315), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT103), .B1(new_n371), .B2(new_n315), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n371), .A2(KEYINPUT103), .A3(new_n315), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n646), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n468), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n551), .B1(new_n558), .B2(new_n559), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n562), .B1(new_n659), .B2(new_n553), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n662), .B(new_n562), .C1(new_n659), .C2(new_n553), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n645), .A2(new_n658), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  AND3_X1   g482(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n449), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT20), .B1(new_n470), .B2(new_n449), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n445), .B1(new_n456), .B2(new_n457), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n437), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n448), .B1(new_n672), .B2(new_n449), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n379), .A3(KEYINPUT104), .A4(new_n469), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n374), .A2(new_n378), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n676), .B1(new_n472), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n645), .A2(new_n665), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NAND2_X1  g496(.A1(new_n295), .A2(new_n296), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n641), .B1(new_n683), .B2(new_n311), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n297), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n582), .A2(KEYINPUT36), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n578), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n593), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n590), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n636), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n565), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  AOI22_X1  g508(.A1(new_n297), .A2(KEYINPUT32), .B1(G472), .B2(new_n312), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n664), .B1(new_n695), .B2(new_n294), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n691), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT105), .B(G900), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n463), .B1(new_n466), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n646), .A2(new_n677), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XNOR2_X1  g517(.A(new_n700), .B(KEYINPUT39), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n643), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n562), .B1(new_n706), .B2(KEYINPUT40), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(KEYINPUT40), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n307), .A2(new_n265), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n302), .A2(new_n267), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n449), .B1(new_n712), .B2(new_n265), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n294), .A2(new_n298), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n689), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT38), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n561), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n379), .A2(new_n646), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n708), .A2(new_n717), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G143), .ZN(G45));
  INV_X1    g537(.A(new_n700), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n646), .A2(new_n656), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n697), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT106), .B(G146), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G48));
  OAI21_X1  g542(.A(new_n311), .B1(new_n619), .B2(new_n622), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n730), .A2(new_n635), .A3(new_n623), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n661), .A2(new_n663), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n314), .A2(new_n595), .A3(new_n732), .A4(new_n658), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT41), .B(G113), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT107), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n733), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n314), .A2(new_n595), .A3(new_n732), .A4(new_n679), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AND4_X1   g552(.A1(new_n663), .A2(new_n661), .A3(new_n689), .A4(new_n731), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n314), .A3(new_n473), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NAND2_X1  g555(.A1(new_n590), .A2(new_n594), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n304), .A2(new_n265), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n188), .B1(new_n743), .B2(new_n288), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n684), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n469), .A3(new_n721), .A4(new_n732), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  INV_X1    g561(.A(new_n725), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n311), .B1(new_n282), .B2(new_n291), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n744), .B1(new_n750), .B2(G472), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n751), .B2(new_n689), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n304), .A2(new_n265), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n189), .B1(new_n753), .B2(new_n271), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n689), .B(new_n754), .C1(new_n640), .C2(new_n641), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n748), .B(new_n732), .C1(new_n752), .C2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT109), .B(G125), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G27));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n297), .B2(KEYINPUT32), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n292), .A2(KEYINPUT110), .A3(new_n293), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n695), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n553), .A3(new_n563), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n643), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n725), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n595), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT42), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n742), .B1(new_n695), .B2(new_n294), .ZN(new_n770));
  INV_X1    g584(.A(new_n766), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n208), .ZN(G33));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n701), .A3(new_n771), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  NAND4_X1  g591(.A1(new_n656), .A2(new_n461), .A3(new_n452), .A4(new_n471), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n779), .A3(KEYINPUT43), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(KEYINPUT44), .A3(new_n642), .A4(new_n689), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n783), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n642), .A2(new_n689), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n765), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n627), .A2(new_n630), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n627), .A2(new_n630), .A3(KEYINPUT45), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n632), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n632), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n801), .A2(new_n623), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n635), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n704), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n785), .A2(KEYINPUT113), .A3(new_n765), .A4(new_n789), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n792), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n635), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n725), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n314), .A2(new_n595), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n765), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  NAND2_X1  g630(.A1(new_n730), .A2(new_n623), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT114), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n811), .B(new_n812), .C1(new_n635), .C2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n782), .A2(new_n463), .A3(new_n783), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n751), .A2(new_n595), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n765), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n716), .A2(new_n595), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n731), .A2(new_n765), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n463), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n824), .A2(new_n656), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n751), .A2(new_n749), .A3(new_n689), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n820), .A2(new_n825), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n828), .A2(new_n674), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n731), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n719), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n822), .A2(new_n563), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n822), .A2(KEYINPUT50), .A3(new_n563), .A4(new_n835), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n823), .B(new_n833), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n256), .A2(G952), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n822), .B2(new_n732), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n784), .A2(new_n463), .A3(new_n826), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n763), .A2(new_n595), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n832), .A2(new_n851), .A3(new_n595), .A4(new_n763), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT48), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n845), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n696), .B(new_n691), .C1(new_n701), .C2(new_n748), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n664), .A2(new_n636), .A3(new_n720), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n690), .A3(new_n724), .A4(new_n715), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n757), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n757), .A2(new_n859), .A3(KEYINPUT52), .A4(new_n861), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n769), .A2(new_n773), .A3(new_n776), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n746), .A2(new_n733), .A3(new_n737), .A4(new_n740), .ZN(new_n868));
  INV_X1    g682(.A(new_n657), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n561), .A2(new_n563), .A3(new_n468), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n645), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n596), .B2(new_n636), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n725), .B1(new_n829), .B2(new_n830), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n377), .A2(new_n372), .A3(new_n700), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n314), .A2(new_n674), .A3(new_n689), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n771), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n742), .A2(new_n636), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n646), .B1(new_n369), .B2(new_n373), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n685), .A2(new_n878), .A3(new_n870), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n692), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n692), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n867), .A2(new_n873), .A3(new_n877), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n858), .B1(new_n866), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n873), .A2(new_n885), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n877), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n769), .A2(new_n773), .A3(new_n776), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n864), .A2(new_n865), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n889), .A2(new_n892), .A3(new_n893), .A4(KEYINPUT53), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n887), .A2(new_n894), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n838), .A2(new_n840), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n833), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n833), .A3(KEYINPUT117), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(KEYINPUT51), .A3(new_n823), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n857), .A2(new_n896), .A3(new_n898), .A4(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n824), .A2(new_n657), .A3(new_n827), .ZN(new_n906));
  OAI22_X1  g720(.A1(new_n905), .A2(new_n906), .B1(G952), .B2(G953), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n818), .B(KEYINPUT49), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n674), .A2(new_n635), .A3(new_n656), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n719), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n595), .A3(new_n562), .A4(new_n716), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n556), .A2(new_n557), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n524), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n311), .B1(new_n887), .B2(new_n894), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n552), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n383), .A2(G952), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n916), .B2(new_n555), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(G51));
  AND3_X1   g737(.A1(new_n887), .A2(new_n895), .A3(new_n894), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n895), .B1(new_n887), .B2(new_n894), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n632), .B(KEYINPUT57), .ZN(new_n927));
  OAI22_X1  g741(.A1(new_n926), .A2(new_n927), .B1(new_n622), .B2(new_n619), .ZN(new_n928));
  INV_X1    g742(.A(new_n798), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n920), .B1(new_n928), .B2(new_n930), .ZN(G54));
  NAND3_X1  g745(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n932), .A2(new_n437), .A3(new_n446), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n437), .B2(new_n446), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n920), .ZN(G60));
  XNOR2_X1  g749(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n315), .A2(new_n449), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n924), .B2(new_n925), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n648), .A2(new_n651), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n920), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n938), .C1(new_n924), .C2(new_n925), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n898), .A2(new_n896), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n945), .A2(new_n946), .A3(new_n942), .A4(new_n938), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n941), .A2(new_n944), .A3(new_n947), .ZN(G63));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT122), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n897), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n591), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n920), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n687), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n949), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n897), .A2(new_n687), .A3(new_n953), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n956), .A2(KEYINPUT61), .A3(new_n957), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(G66));
  NAND2_X1  g778(.A1(new_n888), .A2(new_n383), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  INV_X1    g780(.A(G224), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n467), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n520), .B(new_n523), .C1(G898), .C2(new_n383), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  OAI21_X1  g785(.A(new_n246), .B1(new_n251), .B2(KEYINPUT30), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n441), .Z(new_n973));
  OAI21_X1  g787(.A(G900), .B1(new_n973), .B2(G227), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n464), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n879), .A2(new_n869), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n770), .A2(new_n705), .A3(new_n977), .A4(new_n771), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT124), .Z(new_n979));
  AND2_X1   g793(.A1(new_n757), .A2(new_n859), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n722), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(KEYINPUT62), .A3(new_n722), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n808), .A2(new_n815), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n464), .B(new_n973), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n664), .A2(new_n720), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n805), .A2(new_n849), .A3(new_n704), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n891), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n808), .A2(new_n991), .A3(new_n980), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n808), .B2(new_n980), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n815), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n383), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n987), .B1(new_n995), .B2(new_n973), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n383), .B1(G227), .B2(G900), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT125), .Z(new_n998));
  OAI21_X1  g812(.A(new_n975), .B1(new_n996), .B2(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n994), .B2(new_n888), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n307), .A2(new_n265), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n920), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n985), .A2(new_n986), .A3(new_n889), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n710), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n709), .A2(new_n1001), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1003), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n897), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT127), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n897), .A2(new_n1012), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1004), .A2(new_n1007), .A3(new_n1014), .ZN(G57));
endmodule


