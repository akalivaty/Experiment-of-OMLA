//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1201,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(new_n206), .A2(G50), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n209), .A2(new_n212), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n221), .B(new_n226), .C1(G58), .C2(G232), .ZN(new_n227));
  INV_X1    g0027(.A(new_n214), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT1), .Z(new_n230));
  AOI211_X1 g0030(.A(new_n217), .B(new_n230), .C1(new_n213), .C2(new_n216), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n220), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n201), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n219), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G226), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(G232), .A3(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(G1), .B(G13), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G238), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(KEYINPUT67), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT73), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n266), .B2(new_n271), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT13), .B1(new_n265), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n255), .A2(new_n259), .B1(G238), .B2(new_n263), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT74), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n276), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n277), .A2(KEYINPUT74), .A3(new_n279), .A4(new_n278), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G169), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT14), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n276), .A2(new_n280), .A3(G179), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT14), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n282), .A2(new_n287), .A3(G169), .A4(new_n283), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(G77), .B1(new_n293), .B2(G50), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n290), .B2(G68), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n210), .B1(new_n214), .B2(new_n256), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT11), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n268), .A2(G20), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT69), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n302), .A2(new_n268), .A3(G13), .A4(G20), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n202), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT12), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n303), .ZN(new_n307));
  INV_X1    g0107(.A(new_n296), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n307), .A2(new_n308), .A3(new_n299), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n297), .A2(KEYINPUT11), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n298), .A2(new_n306), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n289), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n250), .A2(G1698), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n314), .B1(new_n246), .B2(new_n250), .C1(new_n315), .C2(new_n223), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n259), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n266), .A2(new_n271), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n263), .A2(G244), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT8), .B(G58), .Z(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n293), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n324), .A2(new_n325), .B1(new_n291), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n290), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n296), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n309), .A2(G77), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n304), .A2(new_n328), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT70), .B(G179), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n322), .B(new_n333), .C1(new_n320), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n320), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT71), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n320), .A2(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n333), .A2(new_n339), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(new_n340), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n313), .A2(new_n336), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n263), .A2(G226), .ZN(new_n346));
  OR2_X1    g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(G1698), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n349), .A2(G222), .B1(new_n352), .B2(G77), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n251), .B1(new_n347), .B2(new_n348), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G223), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n318), .B(new_n346), .C1(new_n356), .C2(new_n258), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n337), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT68), .A2(G58), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT8), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n292), .ZN(new_n362));
  INV_X1    g0162(.A(G150), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n359), .B(new_n362), .C1(new_n363), .C2(new_n325), .ZN(new_n364));
  INV_X1    g0164(.A(G50), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n364), .A2(new_n296), .B1(new_n365), .B2(new_n304), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n309), .A2(G50), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT9), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n345), .A2(new_n358), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT72), .B1(new_n357), .B2(G200), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n370), .B1(new_n369), .B2(new_n368), .C1(new_n358), .C2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(new_n321), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n368), .B(new_n374), .C1(new_n335), .C2(new_n357), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n307), .A2(new_n361), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n352), .B2(new_n290), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n350), .A2(new_n351), .A3(new_n380), .A4(G20), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n293), .A2(G159), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n382), .A2(new_n388), .A3(new_n383), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n390), .B2(new_n296), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n309), .A2(new_n361), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n263), .A2(G232), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n354), .A2(G226), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n349), .A2(G223), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n318), .B(new_n394), .C1(new_n398), .C2(new_n258), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G200), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n399), .A2(new_n337), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n391), .A2(new_n393), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n403));
  NAND2_X1  g0203(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n380), .B1(new_n250), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n352), .A2(KEYINPUT7), .A3(new_n290), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(G68), .B1(G20), .B2(new_n384), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n388), .B1(new_n409), .B2(new_n383), .ZN(new_n410));
  INV_X1    g0210(.A(new_n389), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n296), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n378), .ZN(new_n413));
  AND4_X1   g0213(.A1(new_n412), .A2(new_n401), .A3(new_n413), .A4(new_n393), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT75), .A3(KEYINPUT17), .A4(new_n400), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n399), .A2(new_n321), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n391), .B2(new_n393), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n399), .A2(new_n335), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT18), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n413), .A3(new_n393), .ZN(new_n421));
  AND4_X1   g0221(.A1(KEYINPUT18), .A2(new_n421), .A3(new_n416), .A4(new_n419), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n405), .B(new_n415), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n282), .A2(G200), .A3(new_n283), .ZN(new_n425));
  INV_X1    g0225(.A(new_n312), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n276), .A2(new_n280), .A3(G190), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND4_X1   g0228(.A1(new_n344), .A2(new_n377), .A3(new_n424), .A4(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(G264), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT79), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT79), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n250), .A2(new_n432), .A3(G264), .A4(G1698), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n250), .A2(G257), .A3(new_n251), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n352), .A2(G303), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT80), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n349), .A2(G257), .B1(new_n352), .B2(G303), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT80), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n431), .A4(new_n433), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n259), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n268), .B(G45), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(new_n258), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n268), .A2(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n270), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n446), .A2(G270), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G200), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(G190), .A3(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n304), .A2(new_n219), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n268), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n307), .A2(new_n308), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(G33), .B2(G283), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G33), .B2(new_n224), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n296), .C1(new_n290), .C2(G116), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(new_n460), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n454), .B1(new_n456), .B2(new_n219), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n452), .A2(new_n453), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n321), .B1(new_n442), .B2(new_n450), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT21), .B1(new_n466), .B2(new_n463), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT21), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n468), .B(new_n321), .C1(new_n442), .C2(new_n450), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n442), .A2(G179), .A3(new_n450), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n463), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n451), .A2(KEYINPUT21), .A3(G169), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n470), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n463), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n467), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n290), .B(G87), .C1(new_n350), .C2(new_n351), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n250), .A2(KEYINPUT82), .A3(new_n290), .A4(G87), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT22), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n479), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n481), .A2(new_n482), .A3(new_n486), .A4(KEYINPUT22), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n256), .A2(new_n219), .A3(G20), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT23), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n290), .B2(G107), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n246), .A2(KEYINPUT23), .A3(G20), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(KEYINPUT24), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n296), .A3(new_n500), .ZN(new_n501));
  XOR2_X1   g0301(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n502));
  OR3_X1    g0302(.A1(new_n307), .A2(G107), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n307), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(new_n456), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n349), .A2(G250), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI221_X1 g0309(.A(new_n508), .B1(new_n256), .B2(new_n509), .C1(new_n225), .C2(new_n315), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n259), .B1(G264), .B2(new_n446), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n447), .A2(new_n449), .ZN(new_n512));
  AOI211_X1 g0312(.A(KEYINPUT86), .B(new_n321), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n259), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n446), .A2(G264), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(G169), .ZN(new_n518));
  INV_X1    g0318(.A(G179), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n513), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n507), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n478), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G200), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(G190), .B2(new_n517), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n501), .A2(new_n506), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n445), .A2(G257), .A3(new_n258), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n512), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT77), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT77), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n532), .A3(new_n512), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n354), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n349), .A2(KEYINPUT76), .A3(KEYINPUT4), .A4(G244), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(new_n251), .C1(new_n350), .C2(new_n351), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT76), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n534), .A2(new_n535), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n531), .A2(new_n533), .B1(new_n541), .B2(new_n259), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT78), .B1(new_n542), .B2(new_n525), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n304), .A2(new_n224), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n456), .A2(new_n224), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n246), .B1(new_n406), .B2(new_n407), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n325), .A2(new_n328), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n224), .A2(new_n246), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n246), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n290), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n544), .B(new_n546), .C1(new_n555), .C2(new_n308), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n531), .A2(new_n533), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n541), .A2(new_n259), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT78), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(G200), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n542), .A2(G190), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n543), .A2(new_n557), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(new_n321), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n559), .A3(new_n334), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n556), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n290), .B1(new_n254), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n551), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n290), .B(G68), .C1(new_n350), .C2(new_n351), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n568), .B1(new_n291), .B2(new_n224), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n296), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n304), .A2(new_n326), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n456), .C2(new_n326), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n350), .C2(new_n351), .ZN(new_n579));
  OAI211_X1 g0379(.A(G238), .B(new_n251), .C1(new_n350), .C2(new_n351), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n256), .C2(new_n219), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n259), .ZN(new_n582));
  INV_X1    g0382(.A(new_n449), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n258), .A2(G250), .A3(new_n448), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n334), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n584), .ZN(new_n586));
  AOI211_X1 g0386(.A(new_n449), .B(new_n586), .C1(new_n581), .C2(new_n259), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n578), .B(new_n585), .C1(new_n587), .C2(G169), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n307), .A2(new_n308), .A3(G87), .A4(new_n455), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n576), .A2(new_n577), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n582), .A2(G190), .A3(new_n583), .A4(new_n584), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n587), .C2(new_n525), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n564), .A2(new_n567), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n528), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n524), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n429), .A2(new_n465), .A3(new_n596), .ZN(G372));
  INV_X1    g0397(.A(new_n428), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n415), .A2(new_n405), .ZN(new_n599));
  AOI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n313), .C2(new_n336), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n420), .A2(new_n422), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n373), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n602), .A2(new_n375), .ZN(new_n603));
  INV_X1    g0403(.A(new_n429), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n588), .A2(new_n592), .A3(new_n556), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n565), .A2(new_n566), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT26), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n588), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n588), .A2(new_n592), .A3(new_n556), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n558), .A2(new_n559), .A3(new_n334), .ZN(new_n610));
  AOI21_X1  g0410(.A(G169), .B1(new_n558), .B2(new_n559), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT87), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n565), .A2(new_n613), .A3(new_n566), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n609), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n467), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n472), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n507), .B2(new_n522), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n607), .B(new_n617), .C1(new_n620), .C2(new_n595), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n603), .B1(new_n604), .B2(new_n622), .ZN(G369));
  AOI21_X1  g0423(.A(new_n476), .B1(new_n475), .B2(new_n463), .ZN(new_n624));
  AOI211_X1 g0424(.A(KEYINPUT81), .B(new_n464), .C1(new_n474), .C2(new_n470), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n300), .A2(G20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n268), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n628), .B(KEYINPUT88), .Z(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(G213), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n507), .B1(new_n522), .B2(new_n634), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n528), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT89), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n521), .B1(new_n501), .B2(new_n506), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT90), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n636), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n523), .A2(new_n634), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n645), .ZN(new_n649));
  AOI211_X1 g0449(.A(new_n464), .B(new_n635), .C1(new_n472), .C2(new_n618), .ZN(new_n650));
  INV_X1    g0450(.A(new_n465), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n463), .B2(new_n634), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n478), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n648), .A2(new_n656), .ZN(G399));
  INV_X1    g0457(.A(new_n215), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G41), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n571), .A2(G116), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n209), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT94), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n594), .B(new_n528), .C1(new_n626), .C2(new_n643), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n609), .A2(KEYINPUT26), .A3(new_n612), .A4(new_n614), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n616), .B1(new_n605), .B2(new_n606), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(KEYINPUT93), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n612), .A2(new_n614), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT93), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT26), .A4(new_n609), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n669), .A2(new_n672), .A3(new_n588), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n665), .B1(new_n674), .B2(new_n635), .ZN(new_n675));
  AOI211_X1 g0475(.A(KEYINPUT94), .B(new_n634), .C1(new_n666), .C2(new_n673), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT29), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT95), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT95), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n679), .B(KEYINPUT29), .C1(new_n675), .C2(new_n676), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n621), .A2(new_n635), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT92), .B1(new_n684), .B2(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  NOR4_X1   g0490(.A1(new_n524), .A2(new_n651), .A3(new_n595), .A4(new_n634), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n442), .A2(G179), .A3(new_n450), .A4(new_n587), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n542), .A2(new_n511), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT30), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n542), .A2(new_n335), .A3(new_n587), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n451), .A3(new_n517), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n692), .B2(new_n693), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT31), .B1(new_n700), .B2(new_n634), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT91), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n634), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n691), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n654), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n690), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n664), .B1(new_n715), .B2(G1), .ZN(G364));
  NAND2_X1  g0516(.A1(new_n627), .A2(G45), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n660), .A2(G1), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n290), .A2(G190), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n519), .A3(new_n525), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G159), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT97), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT32), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n290), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n335), .A2(new_n525), .A3(new_n719), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n250), .B1(new_n224), .B2(new_n729), .C1(new_n730), .C2(new_n328), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n525), .A2(G179), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT98), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n290), .A2(new_n337), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n570), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n335), .A2(G20), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n337), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(G50), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n202), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n335), .A2(new_n525), .A3(new_n734), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n731), .B(new_n742), .C1(G58), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n733), .A2(new_n719), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT99), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT99), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G107), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n727), .A2(new_n745), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT100), .Z(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n352), .B1(new_n509), .B2(new_n729), .C1(new_n730), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n740), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n735), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G303), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n724), .A2(G329), .B1(new_n738), .B2(G326), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n761), .B1(new_n762), .B2(new_n749), .C1(new_n763), .C2(new_n743), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n753), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n210), .B1(G20), .B2(new_n321), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n718), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n243), .A2(G45), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n658), .A2(new_n250), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n769), .C1(G45), .C2(new_n209), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n250), .A2(G355), .A3(new_n215), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(G116), .C2(new_n215), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n766), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n775), .B(KEYINPUT101), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n653), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n767), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n718), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n655), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n653), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(G330), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n634), .A2(new_n333), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n343), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n336), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n336), .A2(new_n634), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n621), .A2(new_n635), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n791), .B(KEYINPUT104), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n684), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n712), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n718), .ZN(new_n797));
  INV_X1    g0597(.A(new_n730), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n738), .A2(G303), .B1(new_n798), .B2(G116), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n762), .B2(new_n741), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT102), .Z(new_n801));
  OAI221_X1 g0601(.A(new_n352), .B1(new_n224), .B2(new_n729), .C1(new_n723), .C2(new_n754), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n749), .A2(new_n570), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n735), .A2(new_n246), .B1(new_n743), .B2(new_n509), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT103), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G137), .A2(new_n738), .B1(new_n740), .B2(G150), .ZN(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n743), .C1(new_n809), .C2(new_n730), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT34), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n750), .A2(G68), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n250), .B1(new_n723), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G50), .B2(new_n758), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n729), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n812), .B(new_n818), .C1(G58), .C2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n766), .B1(new_n806), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n821), .A2(new_n781), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n766), .A2(new_n773), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(G77), .B2(new_n824), .C1(new_n774), .C2(new_n792), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n797), .A2(new_n825), .ZN(G384));
  NAND4_X1  g0626(.A1(new_n678), .A2(new_n429), .A3(new_n689), .A4(new_n680), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n603), .ZN(new_n828));
  INV_X1    g0628(.A(new_n632), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n421), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n601), .B2(new_n599), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n421), .A2(new_n416), .A3(new_n419), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n833), .A2(new_n402), .A3(new_n830), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n832), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n837), .B1(new_n423), .B2(new_n831), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(KEYINPUT106), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT39), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n313), .A2(new_n634), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n841), .A2(KEYINPUT106), .A3(KEYINPUT39), .A4(new_n843), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n601), .A2(new_n632), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n841), .A2(new_n843), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n635), .A2(new_n426), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n313), .A2(new_n428), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n312), .B(new_n634), .C1(new_n289), .C2(new_n598), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n793), .A2(new_n790), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n851), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n849), .A2(new_n850), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n828), .B(new_n859), .Z(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n842), .B2(new_n836), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n701), .A2(new_n702), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n792), .B(new_n856), .C1(new_n691), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n861), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n856), .A2(new_n792), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n596), .A2(new_n465), .A3(new_n635), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(new_n865), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(new_n851), .A3(KEYINPUT40), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n865), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n429), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n873), .B(new_n875), .Z(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(G330), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n860), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n268), .B2(new_n627), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n552), .A2(new_n553), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT35), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n212), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n882), .B(G116), .C1(new_n881), .C2(new_n880), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT105), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT36), .ZN(new_n885));
  OAI21_X1  g0685(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n209), .A2(new_n886), .B1(G50), .B2(new_n202), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(G1), .A3(new_n300), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n879), .A2(new_n885), .A3(new_n888), .ZN(G367));
  XOR2_X1   g0689(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n890));
  XOR2_X1   g0690(.A(new_n659), .B(new_n890), .Z(new_n891));
  AND3_X1   g0691(.A1(new_n642), .A2(new_n645), .A3(new_n636), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n646), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT112), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n655), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n655), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n892), .B2(new_n646), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n690), .A2(new_n713), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n670), .A2(new_n556), .A3(new_n634), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT107), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n564), .B(new_n567), .C1(new_n557), .C2(new_n635), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(KEYINPUT107), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n646), .A2(new_n647), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT45), .ZN(new_n909));
  NOR2_X1   g0709(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n648), .B2(new_n906), .ZN(new_n911));
  NAND2_X1  g0711(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n907), .B1(KEYINPUT111), .B2(KEYINPUT44), .C1(new_n646), .C2(new_n647), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(KEYINPUT113), .A3(new_n656), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n656), .A2(KEYINPUT113), .ZN(new_n917));
  INV_X1    g0717(.A(new_n656), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT113), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n909), .A2(new_n914), .A3(new_n917), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n901), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n891), .B1(new_n922), .B2(new_n714), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n717), .A2(G1), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n635), .A2(new_n588), .A3(new_n590), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n593), .B1(new_n635), .B2(new_n590), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT109), .Z(new_n931));
  INV_X1    g0731(.A(KEYINPUT42), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n646), .B2(new_n906), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT108), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n906), .A2(new_n643), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n634), .B1(new_n936), .B2(new_n567), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n646), .A2(new_n932), .A3(new_n906), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT108), .B1(new_n933), .B2(new_n937), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n931), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n931), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(new_n918), .A3(new_n906), .A4(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n948), .A2(new_n944), .B1(new_n656), .B2(new_n907), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n926), .A2(new_n950), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n250), .B1(new_n202), .B2(new_n729), .C1(new_n730), .C2(new_n365), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n741), .A2(new_n809), .B1(new_n363), .B2(new_n743), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G143), .C2(new_n738), .ZN(new_n954));
  INV_X1    g0754(.A(G137), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n723), .A2(new_n955), .B1(new_n735), .B2(new_n201), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT114), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n750), .A2(G77), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(G303), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n352), .B1(new_n246), .B2(new_n729), .C1(new_n743), .C2(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n741), .A2(new_n509), .B1(new_n762), .B2(new_n730), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(G317), .C2(new_n724), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n750), .A2(G97), .ZN(new_n964));
  INV_X1    g0764(.A(new_n738), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n963), .B(new_n964), .C1(new_n754), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n735), .A2(new_n219), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n959), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n766), .ZN(new_n971));
  INV_X1    g0771(.A(new_n769), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n776), .B1(new_n215), .B2(new_n326), .C1(new_n238), .C2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n927), .A2(new_n778), .A3(new_n928), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n971), .A2(new_n781), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n951), .A2(new_n975), .ZN(G387));
  NAND2_X1  g0776(.A1(new_n714), .A2(new_n899), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n659), .A3(new_n901), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n365), .A2(new_n743), .B1(new_n730), .B2(new_n202), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n729), .A2(new_n326), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n250), .B(new_n980), .C1(new_n965), .C2(new_n809), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n979), .B(new_n981), .C1(new_n361), .C2(new_n740), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n723), .A2(new_n363), .B1(new_n735), .B2(new_n328), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT115), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n964), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G303), .A2(new_n798), .B1(new_n744), .B2(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n965), .B2(new_n763), .C1(new_n754), .C2(new_n741), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n762), .B2(new_n729), .C1(new_n509), .C2(new_n735), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n724), .A2(G326), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n352), .B(new_n993), .C1(new_n749), .C2(new_n219), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT116), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n994), .A2(new_n995), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n985), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n323), .A2(new_n365), .ZN(new_n1000));
  AOI211_X1 g0800(.A(G116), .B(new_n571), .C1(new_n1000), .C2(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(G68), .A2(G77), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1001), .A2(new_n261), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n972), .B1(new_n235), .B2(G45), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n661), .A2(new_n352), .A3(new_n658), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(G107), .B2(new_n215), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n999), .A2(new_n766), .B1(new_n776), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n778), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n781), .C1(new_n649), .C2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n899), .B2(new_n925), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n978), .A2(new_n1013), .ZN(G393));
  AOI21_X1  g0814(.A(new_n925), .B1(new_n916), .B2(new_n921), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n907), .A2(new_n775), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n248), .A2(new_n769), .B1(G97), .B2(new_n658), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n776), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n738), .A2(G317), .B1(new_n744), .B2(G311), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT52), .Z(new_n1020));
  OAI21_X1  g0820(.A(new_n352), .B1(new_n735), .B2(new_n762), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n723), .A2(new_n763), .B1(new_n509), .B2(new_n730), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G116), .C2(new_n819), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n740), .A2(G303), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1023), .A3(new_n751), .A4(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n735), .A2(new_n202), .B1(new_n730), .B2(new_n324), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n250), .B1(new_n328), .B2(new_n729), .C1(new_n723), .C2(new_n808), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G50), .C2(new_n740), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n570), .B2(new_n749), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n738), .A2(G150), .B1(new_n744), .B2(G159), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1025), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n718), .B1(new_n1032), .B2(new_n766), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1016), .A2(new_n1018), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT117), .B1(new_n1015), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n919), .B(new_n918), .C1(new_n909), .C2(new_n914), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n921), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n924), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT117), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1034), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n916), .A2(new_n901), .A3(new_n921), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(new_n659), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n715), .B(new_n900), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1042), .A2(new_n1046), .ZN(G390));
  NAND3_X1  g0847(.A1(new_n429), .A2(G330), .A3(new_n874), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n827), .A2(new_n603), .A3(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(G330), .B(new_n792), .C1(new_n691), .C2(new_n710), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT119), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n856), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n871), .A2(G330), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n857), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n712), .A2(new_n792), .A3(new_n856), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n669), .A2(new_n672), .A3(new_n588), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n595), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1059), .B1(new_n524), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT94), .B1(new_n1061), .B2(new_n634), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n674), .A2(new_n665), .A3(new_n635), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n790), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n789), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n854), .A2(KEYINPUT118), .A3(new_n855), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT118), .B1(new_n854), .B2(new_n855), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n874), .A2(G330), .A3(new_n794), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1058), .B(new_n1065), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1057), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1049), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1054), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n846), .A2(new_n848), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n857), .A2(new_n856), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n847), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1064), .A2(new_n789), .A3(new_n1068), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n864), .A2(new_n847), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1073), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n846), .A2(new_n848), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n1058), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1072), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1049), .B(new_n1071), .C1(new_n1086), .C2(new_n1082), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n659), .A3(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n246), .A2(new_n741), .B1(new_n965), .B2(new_n762), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n736), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n250), .B1(new_n819), .B2(G77), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n224), .A2(new_n730), .B1(new_n743), .B2(new_n219), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G294), .B2(new_n724), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n814), .A2(new_n1092), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT54), .B(G143), .Z(new_n1097));
  AOI21_X1  g0897(.A(new_n352), .B1(new_n798), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n809), .B2(new_n729), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n741), .A2(new_n955), .B1(new_n1100), .B2(new_n723), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G128), .C2(new_n738), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n365), .B2(new_n749), .C1(new_n815), .C2(new_n743), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n758), .A2(G150), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1096), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n766), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n361), .B2(new_n824), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n718), .B(new_n1108), .C1(new_n1074), .C2(new_n773), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1087), .A2(new_n1083), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n924), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1090), .A2(new_n1111), .ZN(G378));
  NAND3_X1  g0912(.A1(new_n827), .A2(new_n603), .A3(new_n1048), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT120), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1049), .A2(KEYINPUT120), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1089), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n868), .A2(new_n872), .A3(G330), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n859), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n868), .A2(new_n872), .A3(G330), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(new_n850), .A3(new_n858), .A4(new_n849), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n829), .A2(new_n368), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n377), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n376), .A2(new_n368), .A3(new_n829), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT55), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT55), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1124), .A2(new_n1128), .A3(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT56), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1129), .A3(KEYINPUT56), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1122), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1119), .A2(new_n1133), .A3(new_n1121), .A4(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1117), .A2(KEYINPUT57), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n659), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT57), .B1(new_n1117), .B2(new_n1137), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1143), .A3(new_n659), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1137), .A2(new_n924), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G41), .B1(new_n819), .B2(G68), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n965), .B2(new_n219), .C1(new_n224), .C2(new_n741), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n724), .A2(G283), .B1(G107), .B2(new_n744), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n326), .B2(new_n730), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(G77), .C2(new_n758), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n750), .A2(G58), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n352), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT58), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n365), .B1(new_n350), .B2(G41), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G125), .A2(new_n738), .B1(new_n740), .B2(G132), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n744), .A2(G128), .B1(G150), .B2(new_n819), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n955), .C2(new_n730), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n758), .B2(new_n1097), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT59), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G41), .B1(new_n750), .B2(G159), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G33), .B1(new_n724), .B2(G124), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1154), .A2(new_n1155), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n718), .B1(new_n1164), .B2(new_n766), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(G50), .B2(new_n824), .C1(new_n1134), .C2(new_n774), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1146), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1145), .A2(new_n1168), .ZN(G375));
  AND2_X1   g0969(.A1(new_n1057), .A2(new_n1070), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1113), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(new_n1072), .A3(new_n891), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n723), .A2(new_n1173), .B1(new_n735), .B2(new_n809), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n352), .B(new_n1174), .C1(new_n740), .C2(new_n1097), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n965), .A2(new_n815), .B1(new_n363), .B2(new_n730), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G137), .B2(new_n744), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n819), .A2(G50), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1152), .A4(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n980), .B1(new_n960), .B2(new_n723), .C1(new_n965), .C2(new_n509), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n250), .B(new_n1180), .C1(G283), .C2(new_n744), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n758), .A2(G97), .B1(new_n798), .B2(G107), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n958), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n741), .A2(new_n219), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(new_n766), .B1(new_n202), .B2(new_n823), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n781), .B(new_n1186), .C1(new_n1068), .C2(new_n774), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1170), .B2(new_n925), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1172), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT122), .ZN(G381));
  NOR2_X1   g0991(.A1(new_n1167), .A2(G378), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1145), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n978), .A2(new_n785), .A3(new_n1013), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(G381), .A2(new_n1194), .A3(G384), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n947), .A2(new_n949), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n923), .B2(new_n925), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n975), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(G390), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1193), .A2(new_n1195), .A3(new_n1199), .ZN(G407));
  INV_X1    g1000(.A(G213), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1193), .B2(new_n633), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(G407), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1004(.A(KEYINPUT62), .ZN(new_n1205));
  INV_X1    g1005(.A(G378), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1145), .B2(new_n1168), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT60), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1171), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n659), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1170), .A2(KEYINPUT60), .A3(new_n1113), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1072), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1210), .A2(new_n1212), .A3(KEYINPUT124), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1212), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n660), .B1(new_n1171), .B2(new_n1208), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1189), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G384), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT124), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1215), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G384), .A3(new_n1189), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1117), .A2(new_n891), .A3(new_n1137), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1192), .A2(new_n1226), .B1(G213), .B2(new_n633), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1207), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1205), .B1(new_n1229), .B2(KEYINPUT127), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1144), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1143), .B1(new_n1138), .B2(new_n659), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1141), .ZN(new_n1233));
  OAI21_X1  g1033(.A(G378), .B1(new_n1233), .B2(new_n1167), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G384), .B1(new_n1223), .B2(new_n1189), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1219), .B(new_n1188), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1237), .A3(new_n1227), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(KEYINPUT62), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT61), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1234), .A2(new_n1227), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n633), .A2(G213), .A3(G2897), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1235), .A2(new_n1236), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1243), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1242), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1230), .A2(new_n1240), .A3(new_n1241), .A4(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1194), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n785), .B1(new_n978), .B2(new_n1013), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1041), .A2(new_n1036), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n951), .B2(new_n975), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1199), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(G390), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n951), .A2(new_n1252), .A3(new_n975), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1251), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1248), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1257), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1229), .B2(KEYINPUT63), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1234), .A2(KEYINPUT63), .A3(new_n1227), .A4(new_n1237), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1241), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1225), .A2(new_n1243), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1220), .A2(new_n1224), .A3(new_n1245), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT125), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1242), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1259), .B1(new_n1275), .B2(new_n1238), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1229), .B2(KEYINPUT63), .ZN(new_n1277));
  AND4_X1   g1077(.A1(KEYINPUT126), .A2(new_n1276), .A3(new_n1273), .A4(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1260), .B1(new_n1274), .B2(new_n1278), .ZN(G405));
  NOR2_X1   g1079(.A1(new_n1193), .A2(new_n1207), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1225), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1263), .ZN(G402));
endmodule


