

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757;

  NOR2_X1 U367 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U368 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U369 ( .A(n734), .B(KEYINPUT68), .ZN(n412) );
  AND2_X2 U370 ( .A1(n465), .A2(n632), .ZN(n635) );
  NOR2_X2 U371 ( .A1(n669), .A2(n350), .ZN(n543) );
  XNOR2_X2 U372 ( .A(n530), .B(n529), .ZN(n669) );
  XNOR2_X2 U373 ( .A(n431), .B(KEYINPUT110), .ZN(n693) );
  XNOR2_X2 U374 ( .A(n494), .B(n493), .ZN(n757) );
  NOR2_X1 U375 ( .A1(n682), .A2(n368), .ZN(n437) );
  NOR2_X1 U376 ( .A1(G953), .A2(G237), .ZN(n554) );
  NOR2_X1 U377 ( .A1(n692), .A2(n653), .ZN(n600) );
  XNOR2_X1 U378 ( .A(n437), .B(n584), .ZN(n661) );
  AND2_X1 U379 ( .A1(n457), .A2(n456), .ZN(n464) );
  BUF_X1 U380 ( .A(n719), .Z(n723) );
  NOR2_X1 U381 ( .A1(n373), .A2(n488), .ZN(n487) );
  NAND2_X1 U382 ( .A1(n453), .A2(n452), .ZN(n451) );
  NAND2_X1 U383 ( .A1(n598), .A2(n541), .ZN(n542) );
  BUF_X1 U384 ( .A(n598), .Z(n599) );
  BUF_X1 U385 ( .A(n610), .Z(n630) );
  XNOR2_X1 U386 ( .A(n597), .B(n462), .ZN(n673) );
  OR2_X2 U387 ( .A1(n589), .A2(n391), .ZN(n672) );
  XNOR2_X1 U388 ( .A(n513), .B(KEYINPUT87), .ZN(n744) );
  INV_X2 U389 ( .A(G143), .ZN(n511) );
  INV_X1 U390 ( .A(KEYINPUT3), .ZN(n524) );
  INV_X2 U391 ( .A(G953), .ZN(n748) );
  NAND2_X1 U392 ( .A1(n428), .A2(n474), .ZN(n347) );
  NAND2_X1 U393 ( .A1(n346), .A2(KEYINPUT44), .ZN(n348) );
  NAND2_X1 U394 ( .A1(n347), .A2(n348), .ZN(n469) );
  INV_X1 U395 ( .A(n428), .ZN(n346) );
  XNOR2_X2 U396 ( .A(n449), .B(KEYINPUT32), .ZN(n349) );
  XNOR2_X1 U397 ( .A(n542), .B(KEYINPUT0), .ZN(n350) );
  INV_X1 U398 ( .A(n492), .ZN(n351) );
  BUF_X1 U399 ( .A(n710), .Z(n352) );
  XNOR2_X1 U400 ( .A(n449), .B(KEYINPUT32), .ZN(n387) );
  NAND2_X2 U401 ( .A1(n577), .A2(n476), .ZN(n449) );
  XNOR2_X1 U402 ( .A(n455), .B(n363), .ZN(n728) );
  XNOR2_X1 U403 ( .A(n398), .B(n733), .ZN(n710) );
  XNOR2_X2 U404 ( .A(n400), .B(n447), .ZN(n397) );
  XNOR2_X2 U405 ( .A(n574), .B(KEYINPUT22), .ZN(n577) );
  XNOR2_X2 U406 ( .A(n397), .B(n534), .ZN(n733) );
  NAND2_X1 U407 ( .A1(n438), .A2(n450), .ZN(n406) );
  XNOR2_X1 U408 ( .A(n374), .B(KEYINPUT70), .ZN(n373) );
  NOR2_X1 U409 ( .A1(n647), .A2(n427), .ZN(n426) );
  XNOR2_X1 U410 ( .A(n411), .B(G140), .ZN(n513) );
  INV_X1 U411 ( .A(G137), .ZN(n411) );
  OR2_X1 U412 ( .A1(n713), .A2(G902), .ZN(n389) );
  XNOR2_X1 U413 ( .A(n553), .B(n552), .ZN(n579) );
  NOR2_X1 U414 ( .A1(G902), .A2(n721), .ZN(n553) );
  XNOR2_X1 U415 ( .A(n536), .B(n512), .ZN(n527) );
  XNOR2_X1 U416 ( .A(n571), .B(n460), .ZN(n581) );
  XNOR2_X1 U417 ( .A(n570), .B(n461), .ZN(n460) );
  INV_X1 U418 ( .A(G475), .ZN(n461) );
  NAND2_X1 U419 ( .A1(n408), .A2(KEYINPUT96), .ZN(n402) );
  INV_X1 U420 ( .A(n664), .ZN(n488) );
  INV_X1 U421 ( .A(KEYINPUT44), .ZN(n474) );
  NAND2_X1 U422 ( .A1(G234), .A2(G237), .ZN(n532) );
  XOR2_X1 U423 ( .A(G113), .B(G104), .Z(n559) );
  XOR2_X1 U424 ( .A(G122), .B(G107), .Z(n548) );
  XOR2_X1 U425 ( .A(G140), .B(KEYINPUT11), .Z(n556) );
  XNOR2_X1 U426 ( .A(G143), .B(G122), .ZN(n563) );
  XNOR2_X1 U427 ( .A(n458), .B(G146), .ZN(n537) );
  INV_X1 U428 ( .A(G125), .ZN(n458) );
  AND2_X1 U429 ( .A1(n390), .A2(n597), .ZN(n602) );
  INV_X1 U430 ( .A(n672), .ZN(n390) );
  INV_X1 U431 ( .A(KEYINPUT91), .ZN(n433) );
  NOR2_X1 U432 ( .A1(n435), .A2(n678), .ZN(n434) );
  NOR2_X1 U433 ( .A1(n602), .A2(KEYINPUT91), .ZN(n435) );
  OR2_X1 U434 ( .A1(n725), .A2(G902), .ZN(n498) );
  INV_X1 U435 ( .A(KEYINPUT1), .ZN(n462) );
  XNOR2_X1 U436 ( .A(n396), .B(n478), .ZN(n544) );
  INV_X1 U437 ( .A(KEYINPUT8), .ZN(n478) );
  NAND2_X1 U438 ( .A1(n748), .A2(G234), .ZN(n396) );
  XNOR2_X1 U439 ( .A(n444), .B(n508), .ZN(n443) );
  XOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT76), .Z(n508) );
  XNOR2_X1 U441 ( .A(n507), .B(n445), .ZN(n444) );
  XNOR2_X1 U442 ( .A(G119), .B(KEYINPUT23), .ZN(n507) );
  XNOR2_X1 U443 ( .A(G128), .B(G110), .ZN(n506) );
  XNOR2_X1 U444 ( .A(n537), .B(n497), .ZN(n741) );
  INV_X1 U445 ( .A(KEYINPUT10), .ZN(n497) );
  XNOR2_X1 U446 ( .A(n551), .B(n485), .ZN(n484) );
  XNOR2_X1 U447 ( .A(n486), .B(KEYINPUT7), .ZN(n485) );
  INV_X1 U448 ( .A(KEYINPUT103), .ZN(n486) );
  INV_X1 U449 ( .A(n691), .ZN(n452) );
  XNOR2_X1 U450 ( .A(n388), .B(KEYINPUT39), .ZN(n621) );
  XNOR2_X1 U451 ( .A(n596), .B(n386), .ZN(n385) );
  INV_X1 U452 ( .A(KEYINPUT28), .ZN(n386) );
  OR2_X1 U453 ( .A1(n691), .A2(n391), .ZN(n499) );
  XNOR2_X1 U454 ( .A(n527), .B(n471), .ZN(n713) );
  XNOR2_X1 U455 ( .A(n744), .B(n516), .ZN(n517) );
  NAND2_X1 U456 ( .A1(n747), .A2(n358), .ZN(n395) );
  NOR2_X1 U457 ( .A1(n393), .A2(n392), .ZN(n394) );
  AND2_X1 U458 ( .A1(n358), .A2(n351), .ZN(n392) );
  INV_X1 U459 ( .A(KEYINPUT82), .ZN(n427) );
  INV_X1 U460 ( .A(KEYINPUT46), .ZN(n490) );
  XOR2_X1 U461 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n566) );
  XNOR2_X1 U462 ( .A(KEYINPUT12), .B(KEYINPUT97), .ZN(n565) );
  XOR2_X1 U463 ( .A(KEYINPUT101), .B(KEYINPUT99), .Z(n564) );
  XNOR2_X1 U464 ( .A(KEYINPUT65), .B(G131), .ZN(n558) );
  INV_X1 U465 ( .A(KEYINPUT107), .ZN(n371) );
  INV_X1 U466 ( .A(n692), .ZN(n409) );
  INV_X1 U467 ( .A(n685), .ZN(n670) );
  AND2_X1 U468 ( .A1(n756), .A2(n631), .ZN(n632) );
  INV_X1 U469 ( .A(n665), .ZN(n631) );
  XOR2_X1 U470 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n521) );
  XNOR2_X1 U471 ( .A(G137), .B(G113), .ZN(n520) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n519) );
  XNOR2_X1 U473 ( .A(n446), .B(KEYINPUT88), .ZN(n445) );
  INV_X1 U474 ( .A(KEYINPUT89), .ZN(n446) );
  XNOR2_X1 U475 ( .A(n558), .B(G134), .ZN(n742) );
  XNOR2_X1 U476 ( .A(G902), .B(KEYINPUT15), .ZN(n634) );
  XNOR2_X1 U477 ( .A(n415), .B(n535), .ZN(n414) );
  INV_X1 U478 ( .A(KEYINPUT85), .ZN(n535) );
  XNOR2_X1 U479 ( .A(n412), .B(n417), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT86), .ZN(n419) );
  XNOR2_X1 U482 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n635), .B(KEYINPUT79), .ZN(n667) );
  NOR2_X1 U484 ( .A1(G902), .A2(G237), .ZN(n538) );
  NAND2_X1 U485 ( .A1(n689), .A2(n688), .ZN(n431) );
  AND2_X1 U486 ( .A1(n589), .A2(n357), .ZN(n616) );
  INV_X1 U487 ( .A(n559), .ZN(n447) );
  XNOR2_X1 U488 ( .A(n459), .B(n562), .ZN(n715) );
  XNOR2_X1 U489 ( .A(n569), .B(n561), .ZN(n459) );
  XOR2_X1 U490 ( .A(G104), .B(G107), .Z(n515) );
  XNOR2_X1 U491 ( .A(n399), .B(n536), .ZN(n398) );
  XNOR2_X1 U492 ( .A(n416), .B(n413), .ZN(n399) );
  XNOR2_X1 U493 ( .A(n537), .B(n414), .ZN(n413) );
  BUF_X1 U494 ( .A(n667), .Z(n747) );
  NAND2_X1 U495 ( .A1(n586), .A2(n361), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n442), .B(n440), .ZN(n725) );
  XNOR2_X1 U497 ( .A(n441), .B(n741), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n509), .B(n443), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n547), .B(n483), .ZN(n721) );
  XNOR2_X1 U500 ( .A(n549), .B(n484), .ZN(n483) );
  XOR2_X1 U501 ( .A(G134), .B(KEYINPUT9), .Z(n546) );
  XNOR2_X1 U502 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n493) );
  NAND2_X1 U503 ( .A1(n621), .A2(n657), .ZN(n470) );
  INV_X1 U504 ( .A(KEYINPUT35), .ZN(n439) );
  NOR2_X1 U505 ( .A1(n576), .A2(n578), .ZN(n476) );
  OR2_X1 U506 ( .A1(n379), .A2(n377), .ZN(n653) );
  AND2_X1 U507 ( .A1(n575), .A2(n589), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n711), .B(n463), .ZN(n714) );
  XNOR2_X1 U509 ( .A(n480), .B(n479), .ZN(G51) );
  INV_X1 U510 ( .A(KEYINPUT56), .ZN(n479) );
  NAND2_X1 U511 ( .A1(n481), .A2(n456), .ZN(n480) );
  XNOR2_X1 U512 ( .A(n482), .B(n354), .ZN(n481) );
  NOR2_X1 U513 ( .A1(G953), .A2(n708), .ZN(n709) );
  INV_X1 U514 ( .A(KEYINPUT124), .ZN(n706) );
  XNOR2_X1 U515 ( .A(n475), .B(G122), .ZN(G24) );
  AND2_X1 U516 ( .A1(n705), .A2(n704), .ZN(n353) );
  XOR2_X1 U517 ( .A(n352), .B(n366), .Z(n354) );
  AND2_X1 U518 ( .A1(n432), .A2(n434), .ZN(n355) );
  INV_X1 U519 ( .A(n675), .ZN(n391) );
  XNOR2_X1 U520 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n356) );
  AND2_X1 U521 ( .A1(n603), .A2(n675), .ZN(n357) );
  AND2_X1 U522 ( .A1(n353), .A2(n633), .ZN(n358) );
  AND2_X1 U523 ( .A1(G210), .A2(n540), .ZN(n359) );
  NOR2_X1 U524 ( .A1(n385), .A2(n384), .ZN(n360) );
  AND2_X1 U525 ( .A1(n602), .A2(KEYINPUT91), .ZN(n361) );
  NAND2_X1 U526 ( .A1(n355), .A2(n436), .ZN(n438) );
  XNOR2_X1 U527 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n362) );
  XOR2_X1 U528 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n363) );
  XOR2_X1 U529 ( .A(n638), .B(n637), .Z(n364) );
  XOR2_X1 U530 ( .A(n717), .B(n716), .Z(n365) );
  INV_X1 U531 ( .A(KEYINPUT96), .ZN(n450) );
  NOR2_X1 U532 ( .A1(G952), .A2(n748), .ZN(n727) );
  INV_X1 U533 ( .A(n727), .ZN(n456) );
  XNOR2_X1 U534 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n366) );
  OR2_X1 U535 ( .A1(n634), .A2(n633), .ZN(n367) );
  XNOR2_X1 U536 ( .A(n542), .B(KEYINPUT0), .ZN(n368) );
  XNOR2_X1 U537 ( .A(n542), .B(KEYINPUT0), .ZN(n585) );
  XNOR2_X1 U538 ( .A(n369), .B(n370), .ZN(G57) );
  NAND2_X1 U539 ( .A1(n454), .A2(n456), .ZN(n369) );
  XOR2_X1 U540 ( .A(n640), .B(KEYINPUT114), .Z(n370) );
  XNOR2_X1 U541 ( .A(n372), .B(n371), .ZN(n467) );
  NAND2_X1 U542 ( .A1(n410), .A2(n409), .ZN(n372) );
  NAND2_X1 U543 ( .A1(n748), .A2(G224), .ZN(n415) );
  INV_X1 U544 ( .A(n647), .ZN(n422) );
  NAND2_X1 U545 ( .A1(n719), .A2(G210), .ZN(n482) );
  AND2_X1 U546 ( .A1(n668), .A2(n353), .ZN(n393) );
  AND2_X1 U547 ( .A1(n678), .A2(n616), .ZN(n596) );
  OR2_X1 U548 ( .A1(n638), .A2(G902), .ZN(n472) );
  INV_X1 U549 ( .A(n728), .ZN(n492) );
  NAND2_X1 U550 ( .A1(n710), .A2(n634), .ZN(n539) );
  NAND2_X1 U551 ( .A1(n375), .A2(n651), .ZN(n374) );
  XNOR2_X1 U552 ( .A(n600), .B(KEYINPUT47), .ZN(n375) );
  NOR2_X1 U553 ( .A1(n376), .A2(n385), .ZN(n377) );
  NAND2_X1 U554 ( .A1(n599), .A2(n378), .ZN(n376) );
  NOR2_X1 U555 ( .A1(n384), .A2(n383), .ZN(n378) );
  NAND2_X1 U556 ( .A1(n382), .A2(n380), .ZN(n379) );
  NAND2_X1 U557 ( .A1(n381), .A2(n383), .ZN(n380) );
  NAND2_X1 U558 ( .A1(n599), .A2(n597), .ZN(n381) );
  NAND2_X1 U559 ( .A1(n385), .A2(n383), .ZN(n382) );
  INV_X1 U560 ( .A(KEYINPUT77), .ZN(n383) );
  INV_X1 U561 ( .A(n597), .ZN(n384) );
  NAND2_X1 U562 ( .A1(n387), .A2(n422), .ZN(n421) );
  NAND2_X1 U563 ( .A1(n426), .A2(n349), .ZN(n424) );
  XNOR2_X1 U564 ( .A(n349), .B(G119), .ZN(G21) );
  NAND2_X1 U565 ( .A1(n611), .A2(n689), .ZN(n388) );
  XNOR2_X1 U566 ( .A(n606), .B(KEYINPUT74), .ZN(n611) );
  XNOR2_X2 U567 ( .A(n389), .B(G469), .ZN(n597) );
  XNOR2_X2 U568 ( .A(n498), .B(n510), .ZN(n589) );
  NAND2_X1 U569 ( .A1(n394), .A2(n395), .ZN(n707) );
  NAND2_X1 U570 ( .A1(n544), .A2(G221), .ZN(n441) );
  XNOR2_X2 U571 ( .A(G110), .B(KEYINPUT84), .ZN(n734) );
  XNOR2_X1 U572 ( .A(n528), .B(n400), .ZN(n473) );
  XNOR2_X2 U573 ( .A(n526), .B(n356), .ZN(n400) );
  XNOR2_X2 U574 ( .A(n401), .B(KEYINPUT72), .ZN(n583) );
  NOR2_X2 U575 ( .A1(n673), .A2(n672), .ZN(n401) );
  INV_X1 U576 ( .A(n661), .ZN(n407) );
  NAND2_X1 U577 ( .A1(n403), .A2(n402), .ZN(n410) );
  NAND2_X1 U578 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U579 ( .A1(n661), .A2(n450), .ZN(n404) );
  NAND2_X1 U580 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U581 ( .A(n438), .ZN(n408) );
  XNOR2_X1 U582 ( .A(n412), .B(n517), .ZN(n471) );
  XNOR2_X2 U583 ( .A(n420), .B(KEYINPUT19), .ZN(n598) );
  NOR2_X1 U584 ( .A1(n624), .A2(n420), .ZN(n617) );
  NAND2_X2 U585 ( .A1(n610), .A2(n688), .ZN(n420) );
  NAND2_X1 U586 ( .A1(n421), .A2(n427), .ZN(n425) );
  NAND2_X1 U587 ( .A1(n423), .A2(n475), .ZN(n428) );
  NAND2_X1 U588 ( .A1(n425), .A2(n424), .ZN(n423) );
  NAND2_X1 U589 ( .A1(n429), .A2(n430), .ZN(n466) );
  XNOR2_X1 U590 ( .A(n591), .B(KEYINPUT78), .ZN(n429) );
  INV_X1 U591 ( .A(n667), .ZN(n430) );
  NAND2_X1 U592 ( .A1(n612), .A2(n613), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n491), .B(n490), .ZN(n489) );
  NAND2_X1 U594 ( .A1(n350), .A2(n433), .ZN(n432) );
  AND2_X1 U595 ( .A1(n589), .A2(n391), .ZN(n676) );
  XNOR2_X2 U596 ( .A(n573), .B(n439), .ZN(n475) );
  AND2_X1 U597 ( .A1(n577), .A2(n448), .ZN(n647) );
  AND2_X2 U598 ( .A1(n496), .A2(n495), .ZN(n719) );
  NAND2_X1 U599 ( .A1(n719), .A2(G475), .ZN(n718) );
  XNOR2_X2 U600 ( .A(n451), .B(KEYINPUT41), .ZN(n685) );
  INV_X1 U601 ( .A(n693), .ZN(n453) );
  XNOR2_X1 U602 ( .A(n639), .B(n364), .ZN(n454) );
  NAND2_X1 U603 ( .A1(n469), .A2(n468), .ZN(n455) );
  XNOR2_X2 U604 ( .A(n630), .B(n609), .ZN(n689) );
  XNOR2_X1 U605 ( .A(n718), .B(n365), .ZN(n457) );
  XNOR2_X1 U606 ( .A(n713), .B(n712), .ZN(n463) );
  XNOR2_X1 U607 ( .A(n464), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U608 ( .A1(n685), .A2(n360), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n619), .B(n620), .ZN(n465) );
  NAND2_X1 U610 ( .A1(n466), .A2(n367), .ZN(n496) );
  AND2_X1 U611 ( .A1(n467), .A2(n590), .ZN(n468) );
  XNOR2_X2 U612 ( .A(G119), .B(G116), .ZN(n525) );
  NOR2_X2 U613 ( .A1(n728), .A2(n634), .ZN(n591) );
  INV_X1 U614 ( .A(n755), .ZN(n613) );
  XNOR2_X2 U615 ( .A(n470), .B(n362), .ZN(n755) );
  XNOR2_X2 U616 ( .A(n472), .B(G472), .ZN(n678) );
  XNOR2_X1 U617 ( .A(n527), .B(n473), .ZN(n638) );
  XNOR2_X2 U618 ( .A(n539), .B(n359), .ZN(n610) );
  NAND2_X1 U619 ( .A1(n577), .A2(n614), .ZN(n477) );
  NOR2_X1 U620 ( .A1(n477), .A2(n625), .ZN(n587) );
  NAND2_X1 U621 ( .A1(n544), .A2(G217), .ZN(n545) );
  XNOR2_X2 U622 ( .A(n745), .B(G101), .ZN(n536) );
  XNOR2_X2 U623 ( .A(n550), .B(KEYINPUT4), .ZN(n745) );
  NAND2_X1 U624 ( .A1(n489), .A2(n487), .ZN(n619) );
  INV_X1 U625 ( .A(n668), .ZN(n495) );
  NOR2_X2 U626 ( .A1(n585), .A2(n499), .ZN(n574) );
  XNOR2_X1 U627 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n742), .B(G146), .ZN(n512) );
  XOR2_X1 U629 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n502) );
  NAND2_X1 U630 ( .A1(n634), .A2(G234), .ZN(n500) );
  XNOR2_X1 U631 ( .A(n500), .B(KEYINPUT20), .ZN(n503) );
  NAND2_X1 U632 ( .A1(n503), .A2(G221), .ZN(n501) );
  XNOR2_X1 U633 ( .A(n502), .B(n501), .ZN(n675) );
  XOR2_X1 U634 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n505) );
  NAND2_X1 U635 ( .A1(n503), .A2(G217), .ZN(n504) );
  XNOR2_X1 U636 ( .A(n505), .B(n504), .ZN(n510) );
  XNOR2_X1 U637 ( .A(n506), .B(n513), .ZN(n509) );
  XNOR2_X2 U638 ( .A(n511), .B(G128), .ZN(n550) );
  NAND2_X1 U639 ( .A1(G227), .A2(n748), .ZN(n514) );
  XNOR2_X1 U640 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U641 ( .A1(n554), .A2(G210), .ZN(n518) );
  XNOR2_X1 U642 ( .A(n519), .B(n518), .ZN(n523) );
  XNOR2_X1 U643 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U644 ( .A(n523), .B(n522), .Z(n528) );
  XOR2_X1 U645 ( .A(n678), .B(KEYINPUT6), .Z(n576) );
  NAND2_X1 U646 ( .A1(n583), .A2(n576), .ZN(n530) );
  AND2_X1 U647 ( .A1(n748), .A2(G952), .ZN(n594) );
  NAND2_X1 U648 ( .A1(G953), .A2(G902), .ZN(n592) );
  NOR2_X1 U649 ( .A1(G898), .A2(n592), .ZN(n531) );
  NOR2_X1 U650 ( .A1(n594), .A2(n531), .ZN(n533) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n532), .Z(n702) );
  NOR2_X1 U652 ( .A1(n533), .A2(n702), .ZN(n541) );
  XOR2_X1 U653 ( .A(n548), .B(KEYINPUT16), .Z(n534) );
  XNOR2_X1 U654 ( .A(n538), .B(KEYINPUT73), .ZN(n540) );
  NAND2_X1 U655 ( .A1(G214), .A2(n540), .ZN(n688) );
  XNOR2_X1 U656 ( .A(n543), .B(KEYINPUT34), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U658 ( .A(G116), .B(n548), .ZN(n549) );
  INV_X1 U659 ( .A(n550), .ZN(n551) );
  XNOR2_X1 U660 ( .A(KEYINPUT104), .B(G478), .ZN(n552) );
  NAND2_X1 U661 ( .A1(G214), .A2(n554), .ZN(n555) );
  XNOR2_X1 U662 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U663 ( .A(n557), .B(n741), .Z(n562) );
  INV_X1 U664 ( .A(n558), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U666 ( .A(n564), .B(n563), .ZN(n568) );
  XNOR2_X1 U667 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U668 ( .A(n568), .B(n567), .Z(n569) );
  NOR2_X1 U669 ( .A1(G902), .A2(n715), .ZN(n571) );
  XNOR2_X1 U670 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n570) );
  NOR2_X1 U671 ( .A1(n579), .A2(n581), .ZN(n607) );
  NAND2_X1 U672 ( .A1(n572), .A2(n607), .ZN(n573) );
  INV_X1 U673 ( .A(n673), .ZN(n625) );
  NOR2_X1 U674 ( .A1(n678), .A2(n625), .ZN(n575) );
  NAND2_X1 U675 ( .A1(n579), .A2(n581), .ZN(n691) );
  NAND2_X1 U676 ( .A1(n589), .A2(n625), .ZN(n578) );
  INV_X1 U677 ( .A(n576), .ZN(n614) );
  INV_X1 U678 ( .A(n579), .ZN(n580) );
  NOR2_X1 U679 ( .A1(n581), .A2(n580), .ZN(n657) );
  NAND2_X1 U680 ( .A1(n581), .A2(n580), .ZN(n648) );
  XNOR2_X1 U681 ( .A(KEYINPUT105), .B(n648), .ZN(n622) );
  NOR2_X1 U682 ( .A1(n657), .A2(n622), .ZN(n582) );
  XNOR2_X1 U683 ( .A(n582), .B(KEYINPUT106), .ZN(n692) );
  NAND2_X1 U684 ( .A1(n678), .A2(n583), .ZN(n682) );
  XNOR2_X1 U685 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n584) );
  INV_X1 U686 ( .A(n368), .ZN(n586) );
  XNOR2_X1 U687 ( .A(n587), .B(KEYINPUT81), .ZN(n588) );
  NOR2_X1 U688 ( .A1(n589), .A2(n588), .ZN(n641) );
  INV_X1 U689 ( .A(n641), .ZN(n590) );
  XOR2_X1 U690 ( .A(KEYINPUT48), .B(KEYINPUT80), .Z(n620) );
  NOR2_X1 U691 ( .A1(G900), .A2(n592), .ZN(n593) );
  NOR2_X1 U692 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U693 ( .A1(n595), .A2(n702), .ZN(n603) );
  NAND2_X1 U694 ( .A1(n678), .A2(n688), .ZN(n601) );
  XNOR2_X1 U695 ( .A(KEYINPUT30), .B(n601), .ZN(n605) );
  NAND2_X1 U696 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U697 ( .A1(n611), .A2(n607), .ZN(n608) );
  NAND2_X1 U698 ( .A1(n630), .A2(n608), .ZN(n651) );
  XNOR2_X1 U699 ( .A(KEYINPUT71), .B(KEYINPUT38), .ZN(n609) );
  INV_X1 U700 ( .A(n757), .ZN(n612) );
  INV_X1 U701 ( .A(n657), .ZN(n654) );
  NOR2_X1 U702 ( .A1(n654), .A2(n614), .ZN(n615) );
  NAND2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n617), .B(KEYINPUT36), .ZN(n618) );
  NAND2_X1 U705 ( .A1(n618), .A2(n625), .ZN(n664) );
  NAND2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U707 ( .A(KEYINPUT112), .B(n623), .ZN(n756) );
  XOR2_X1 U708 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n628) );
  NOR2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n626), .A2(n688), .ZN(n627) );
  XNOR2_X1 U711 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n665) );
  INV_X1 U713 ( .A(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n635), .A2(KEYINPUT2), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n351), .A2(n636), .ZN(n668) );
  NAND2_X1 U716 ( .A1(n719), .A2(G472), .ZN(n639) );
  XOR2_X1 U717 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n637) );
  INV_X1 U718 ( .A(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U719 ( .A(G101), .B(n641), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT115), .ZN(G3) );
  NAND2_X1 U721 ( .A1(n408), .A2(n657), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n643), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n645) );
  INV_X1 U724 ( .A(n648), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n408), .A2(n660), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U727 ( .A(G107), .B(n646), .ZN(G9) );
  XOR2_X1 U728 ( .A(G110), .B(n647), .Z(G12) );
  NOR2_X1 U729 ( .A1(n648), .A2(n653), .ZN(n650) );
  XNOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .ZN(n649) );
  XNOR2_X1 U731 ( .A(n650), .B(n649), .ZN(G30) );
  XNOR2_X1 U732 ( .A(G143), .B(KEYINPUT116), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(G45) );
  NOR2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n656) );
  XNOR2_X1 U735 ( .A(G146), .B(KEYINPUT117), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n656), .B(n655), .ZN(G48) );
  NAND2_X1 U737 ( .A1(n661), .A2(n657), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(KEYINPUT118), .ZN(n659) );
  XNOR2_X1 U739 ( .A(G113), .B(n659), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n662), .B(G116), .ZN(G18) );
  XOR2_X1 U742 ( .A(G125), .B(KEYINPUT37), .Z(n663) );
  XNOR2_X1 U743 ( .A(n664), .B(n663), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G140), .B(n665), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT119), .ZN(G42) );
  NOR2_X1 U746 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U747 ( .A(n671), .B(KEYINPUT123), .ZN(n705) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n674), .ZN(n680) );
  XOR2_X1 U750 ( .A(KEYINPUT49), .B(n676), .Z(n677) );
  NOR2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n681), .B(KEYINPUT120), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n684), .Z(n686) );
  NAND2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U757 ( .A(KEYINPUT121), .B(n687), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U762 ( .A1(n669), .A2(n696), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT122), .ZN(n698) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U765 ( .A(n700), .B(KEYINPUT52), .ZN(n701) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n703), .A2(G952), .ZN(n704) );
  XNOR2_X1 U768 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U769 ( .A(KEYINPUT53), .B(n709), .ZN(G75) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  NAND2_X1 U771 ( .A1(n723), .A2(G469), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n727), .A2(n714), .ZN(G54) );
  XNOR2_X1 U773 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n715), .B(KEYINPUT126), .ZN(n716) );
  NAND2_X1 U775 ( .A1(G478), .A2(n723), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n727), .A2(n722), .ZN(G63) );
  NAND2_X1 U778 ( .A1(G217), .A2(n723), .ZN(n724) );
  XNOR2_X1 U779 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(G66) );
  OR2_X1 U781 ( .A1(G953), .A2(n351), .ZN(n732) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U783 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n733), .B(G101), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n734), .B(n735), .ZN(n737) );
  NOR2_X1 U788 ( .A1(G898), .A2(n748), .ZN(n736) );
  NOR2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U791 ( .A(KEYINPUT127), .B(n740), .Z(G69) );
  XOR2_X1 U792 ( .A(n742), .B(n741), .Z(n743) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n746) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n750) );
  XNOR2_X1 U795 ( .A(n747), .B(n750), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n754) );
  XNOR2_X1 U797 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G953), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U801 ( .A(G131), .B(n755), .Z(G33) );
  XNOR2_X1 U802 ( .A(G134), .B(n756), .ZN(G36) );
  XOR2_X1 U803 ( .A(n757), .B(G137), .Z(G39) );
endmodule

