

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U323 ( .A1(n564), .A2(n561), .ZN(n455) );
  AND2_X1 U324 ( .A1(n518), .A2(n411), .ZN(n568) );
  XOR2_X2 U325 ( .A(n360), .B(n359), .Z(n561) );
  XOR2_X1 U326 ( .A(n309), .B(n308), .Z(n574) );
  XNOR2_X1 U327 ( .A(n379), .B(n378), .ZN(n396) );
  NOR2_X1 U328 ( .A1(n396), .A2(n542), .ZN(n397) );
  NOR2_X1 U329 ( .A1(n545), .A2(n398), .ZN(n399) );
  XNOR2_X1 U330 ( .A(n440), .B(n295), .ZN(n296) );
  XNOR2_X1 U331 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U332 ( .A(n451), .B(G176GAT), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n292) );
  XNOR2_X1 U335 ( .A(KEYINPUT72), .B(KEYINPUT74), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n299) );
  XOR2_X1 U337 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n294) );
  XNOR2_X1 U338 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n297) );
  XOR2_X1 U340 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  AND2_X1 U341 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n309) );
  XNOR2_X1 U343 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n300), .B(KEYINPUT13), .ZN(n383) );
  XOR2_X1 U345 ( .A(KEYINPUT73), .B(G92GAT), .Z(n302) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G85GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n345) );
  XOR2_X1 U348 ( .A(n383), .B(n345), .Z(n307) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n303), .B(G148GAT), .ZN(n421) );
  XOR2_X1 U351 ( .A(G64GAT), .B(KEYINPUT75), .Z(n305) );
  XNOR2_X1 U352 ( .A(G176GAT), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n335) );
  XNOR2_X1 U354 ( .A(n421), .B(n335), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n574), .B(KEYINPUT41), .Z(n537) );
  INV_X1 U357 ( .A(n537), .ZN(n554) );
  XOR2_X1 U358 ( .A(G85GAT), .B(G155GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(G127GAT), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U361 ( .A(G29GAT), .B(G162GAT), .Z(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n327) );
  XOR2_X1 U363 ( .A(G57GAT), .B(KEYINPUT5), .Z(n315) );
  XNOR2_X1 U364 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U366 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n317) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(G148GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U369 ( .A(n319), .B(n318), .Z(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n321) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(G134GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n437) );
  XOR2_X1 U373 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n323) );
  XNOR2_X1 U374 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n418) );
  XNOR2_X1 U376 ( .A(n437), .B(n418), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n329) );
  NAND2_X1 U379 ( .A1(G225GAT), .A2(G233GAT), .ZN(n328) );
  XOR2_X1 U380 ( .A(n329), .B(n328), .Z(n518) );
  XOR2_X1 U381 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n331) );
  NAND2_X1 U382 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(n332), .B(G92GAT), .Z(n337) );
  XOR2_X1 U385 ( .A(G211GAT), .B(KEYINPUT21), .Z(n334) );
  XNOR2_X1 U386 ( .A(G197GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n417) );
  XNOR2_X1 U388 ( .A(n417), .B(n335), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n344) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n338), .B(KEYINPUT79), .ZN(n348) );
  XOR2_X1 U392 ( .A(G183GAT), .B(KEYINPUT80), .Z(n386) );
  XOR2_X1 U393 ( .A(n348), .B(n386), .Z(n342) );
  XOR2_X1 U394 ( .A(G169GAT), .B(G8GAT), .Z(n366) );
  XOR2_X1 U395 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n340) );
  XNOR2_X1 U396 ( .A(KEYINPUT86), .B(KEYINPUT18), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n435) );
  XNOR2_X1 U398 ( .A(n366), .B(n435), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n495) );
  INV_X1 U401 ( .A(n495), .ZN(n522) );
  INV_X1 U402 ( .A(KEYINPUT48), .ZN(n409) );
  XOR2_X1 U403 ( .A(n345), .B(G106GAT), .Z(n347) );
  XOR2_X1 U404 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U405 ( .A(G218GAT), .B(n424), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n352) );
  XOR2_X1 U407 ( .A(n348), .B(KEYINPUT10), .Z(n350) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U410 ( .A(n352), .B(n351), .Z(n360) );
  XOR2_X1 U411 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n354) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(G29GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(KEYINPUT7), .B(n355), .Z(n373) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n357) );
  XNOR2_X1 U416 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n373), .B(n358), .ZN(n359) );
  INV_X1 U419 ( .A(n561), .ZN(n545) );
  XOR2_X1 U420 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n362) );
  XNOR2_X1 U421 ( .A(G197GAT), .B(G1GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n377) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G141GAT), .Z(n364) );
  XNOR2_X1 U424 ( .A(G15GAT), .B(G113GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U426 ( .A(n365), .B(G50GAT), .Z(n368) );
  XNOR2_X1 U427 ( .A(n366), .B(G36GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U429 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n370) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U432 ( .A(n372), .B(n371), .Z(n375) );
  XNOR2_X1 U433 ( .A(n373), .B(KEYINPUT30), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U435 ( .A(n377), .B(n376), .Z(n534) );
  NAND2_X1 U436 ( .A1(n534), .A2(n537), .ZN(n379) );
  XOR2_X1 U437 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n378) );
  XOR2_X1 U438 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n385) );
  XOR2_X1 U439 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n381) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(G64GAT), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U444 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U445 ( .A(n386), .B(n423), .Z(n388) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U448 ( .A(n390), .B(n389), .Z(n395) );
  XOR2_X1 U449 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XOR2_X1 U450 ( .A(G78GAT), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U451 ( .A(G1GAT), .B(G71GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n441), .B(n393), .ZN(n394) );
  XOR2_X1 U454 ( .A(n395), .B(n394), .Z(n578) );
  INV_X1 U455 ( .A(n578), .ZN(n542) );
  XNOR2_X1 U456 ( .A(n397), .B(KEYINPUT115), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(KEYINPUT47), .ZN(n407) );
  XOR2_X1 U458 ( .A(KEYINPUT45), .B(KEYINPUT65), .Z(n402) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n400) );
  XOR2_X1 U460 ( .A(n561), .B(n400), .Z(n581) );
  NAND2_X1 U461 ( .A1(n542), .A2(n581), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n403), .B(KEYINPUT116), .ZN(n404) );
  NOR2_X1 U464 ( .A1(n574), .A2(n404), .ZN(n405) );
  INV_X1 U465 ( .A(n534), .ZN(n569) );
  NAND2_X1 U466 ( .A1(n405), .A2(n569), .ZN(n406) );
  NAND2_X1 U467 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n549) );
  NOR2_X1 U469 ( .A1(n522), .A2(n549), .ZN(n410) );
  XNOR2_X1 U470 ( .A(KEYINPUT54), .B(n410), .ZN(n411) );
  XOR2_X1 U471 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n428) );
  XOR2_X1 U474 ( .A(G204GAT), .B(KEYINPUT22), .Z(n415) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U477 ( .A(n416), .B(KEYINPUT89), .Z(n420) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n472) );
  NAND2_X1 U484 ( .A1(n568), .A2(n472), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n429), .B(KEYINPUT122), .ZN(n430) );
  XNOR2_X1 U486 ( .A(KEYINPUT55), .B(n430), .ZN(n450) );
  XOR2_X1 U487 ( .A(G176GAT), .B(G183GAT), .Z(n432) );
  XNOR2_X1 U488 ( .A(KEYINPUT87), .B(KEYINPUT84), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n449) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n434) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n439) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT64), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G190GAT), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n524) );
  INV_X1 U503 ( .A(n524), .ZN(n532) );
  NAND2_X1 U504 ( .A1(n450), .A2(n532), .ZN(n564) );
  NOR2_X1 U505 ( .A1(n554), .A2(n564), .ZN(n453) );
  XNOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n451) );
  INV_X1 U507 ( .A(G190GAT), .ZN(n457) );
  XNOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  NOR2_X1 U511 ( .A1(n569), .A2(n574), .ZN(n489) );
  XOR2_X1 U512 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n459) );
  NAND2_X1 U513 ( .A1(n542), .A2(n561), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n475) );
  NOR2_X1 U515 ( .A1(n524), .A2(n522), .ZN(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT97), .B(n460), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n461), .A2(n472), .ZN(n464) );
  XNOR2_X1 U518 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n468) );
  NOR2_X1 U521 ( .A1(n472), .A2(n532), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n465), .B(KEYINPUT26), .ZN(n567) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n466) );
  XOR2_X1 U524 ( .A(n466), .B(n495), .Z(n470) );
  NAND2_X1 U525 ( .A1(n567), .A2(n470), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n518), .ZN(n474) );
  INV_X1 U528 ( .A(n518), .ZN(n492) );
  NAND2_X1 U529 ( .A1(n470), .A2(n492), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT96), .ZN(n550) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT28), .ZN(n526) );
  INV_X1 U532 ( .A(n526), .ZN(n499) );
  NOR2_X1 U533 ( .A1(n550), .A2(n499), .ZN(n531) );
  NAND2_X1 U534 ( .A1(n531), .A2(n524), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n486) );
  AND2_X1 U536 ( .A1(n475), .A2(n486), .ZN(n503) );
  NAND2_X1 U537 ( .A1(n489), .A2(n503), .ZN(n482) );
  NOR2_X1 U538 ( .A1(n518), .A2(n482), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n478), .Z(G1324GAT) );
  NOR2_X1 U542 ( .A1(n522), .A2(n482), .ZN(n479) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n524), .A2(n482), .ZN(n481) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U547 ( .A1(n526), .A2(n482), .ZN(n483) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n485) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n485), .B(n484), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n581), .A2(n486), .ZN(n487) );
  NOR2_X1 U553 ( .A1(n542), .A2(n487), .ZN(n488) );
  XOR2_X1 U554 ( .A(KEYINPUT37), .B(n488), .Z(n515) );
  NAND2_X1 U555 ( .A1(n489), .A2(n515), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n490), .B(KEYINPUT38), .ZN(n491) );
  XNOR2_X1 U557 ( .A(KEYINPUT103), .B(n491), .ZN(n500) );
  NAND2_X1 U558 ( .A1(n492), .A2(n500), .ZN(n493) );
  XOR2_X1 U559 ( .A(n494), .B(n493), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n495), .A2(n500), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n500), .A2(n532), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U567 ( .A1(n537), .A2(n569), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n502), .B(KEYINPUT105), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n516), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(KEYINPUT106), .B(n504), .ZN(n512) );
  NOR2_X1 U571 ( .A1(n512), .A2(n518), .ZN(n506) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n512), .A2(n522), .ZN(n508) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(n508), .Z(n509) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n512), .A2(n524), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n510) );
  XNOR2_X1 U580 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n512), .A2(n526), .ZN(n514) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(KEYINPUT110), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n527), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n522), .ZN(n523) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n524), .ZN(n525) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U595 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XOR2_X1 U598 ( .A(G113GAT), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n549), .A2(n533), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n546), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U604 ( .A1(n546), .A2(n537), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT118), .Z(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n546), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n551), .A2(n567), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n569), .A2(n560), .ZN(n552) );
  XOR2_X1 U617 ( .A(KEYINPUT120), .B(n552), .Z(n553) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  NOR2_X1 U619 ( .A1(n560), .A2(n554), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n578), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NOR2_X1 U628 ( .A1(n569), .A2(n564), .ZN(n563) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n563), .Z(G1348GAT) );
  NOR2_X1 U630 ( .A1(n578), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n577) );
  NOR2_X1 U634 ( .A1(n577), .A2(n569), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  INV_X1 U639 ( .A(n577), .ZN(n582) );
  AND2_X1 U640 ( .A1(n574), .A2(n582), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(n579), .Z(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

