//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .A3(G137), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(new_n465), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT65), .B1(new_n469), .B2(new_n470), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n464), .A2(new_n479), .A3(new_n465), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(G125), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n468), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n464), .A2(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n466), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n485), .A2(G126), .A3(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n468), .A2(G138), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n478), .A2(new_n480), .A3(new_n495), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(G88), .A2(new_n517), .B1(new_n518), .B2(G50), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n509), .A2(G62), .ZN(new_n521));
  AND2_X1   g096(.A1(G75), .A2(G543), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n520), .B(G651), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT69), .B1(new_n524), .B2(new_n510), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n517), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n518), .A2(G51), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n509), .A2(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n509), .A2(new_n516), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n516), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n537), .A2(new_n545), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n509), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n517), .B2(G91), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n539), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n516), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G299));
  OR2_X1    g141(.A1(new_n541), .A2(new_n543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT70), .ZN(G301));
  NAND3_X1  g143(.A1(new_n517), .A2(KEYINPUT71), .A3(G87), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n537), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n509), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(G651), .A2(new_n574), .B1(new_n518), .B2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G288));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n537), .A2(new_n577), .B1(new_n539), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n509), .A2(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n510), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(G305));
  XNOR2_X1  g160(.A(KEYINPUT74), .B(G85), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT73), .B(G47), .Z(new_n587));
  OAI22_X1  g162(.A1(new_n537), .A2(new_n586), .B1(new_n539), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n510), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND3_X1  g167(.A1(new_n509), .A2(new_n516), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n557), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n518), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  XNOR2_X1  g176(.A(G171), .B(KEYINPUT70), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G284));
  AOI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G286), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(G299), .B(KEYINPUT75), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(G297));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n605), .ZN(G280));
  INV_X1    g184(.A(new_n600), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(new_n550), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n605), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n600), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n478), .A2(new_n480), .ZN(new_n618));
  NOR3_X1   g193(.A1(new_n618), .A2(new_n463), .A3(G2105), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n487), .A2(G123), .B1(G135), .B2(new_n466), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n629), .A2(new_n468), .A3(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n468), .B2(G111), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n628), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n626), .A2(new_n627), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT77), .Z(G156));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT79), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  AOI21_X1  g216(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  AOI21_X1  g234(.A(new_n657), .B1(new_n656), .B2(KEYINPUT81), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(KEYINPUT81), .B2(new_n656), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n656), .B(KEYINPUT17), .Z(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n655), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n671), .A2(new_n674), .A3(new_n678), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G6), .A2(G16), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n583), .B(KEYINPUT72), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G16), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G22), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT84), .Z(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G303), .B2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(G23), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n573), .A2(new_n575), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n704), .A2(new_n705), .B1(new_n698), .B2(new_n697), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n693), .A2(new_n699), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n693), .A2(new_n709), .A3(new_n699), .A4(new_n706), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n694), .A2(G24), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT83), .Z(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n591), .B2(new_n694), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1986), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n487), .A2(G119), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n466), .A2(G131), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n710), .A2(KEYINPUT85), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(KEYINPUT85), .B1(new_n710), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n708), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(KEYINPUT36), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(new_n708), .C1(new_n728), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n735));
  OR3_X1    g310(.A1(new_n735), .A2(G5), .A3(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(G5), .B2(G16), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n736), .B(new_n737), .C1(new_n567), .C2(new_n694), .ZN(new_n738));
  INV_X1    g313(.A(G1961), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n694), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n694), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT88), .B(G1966), .Z(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n466), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  INV_X1    g322(.A(G129), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n747), .C1(new_n486), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n715), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n715), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n694), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n550), .B2(new_n694), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n756), .A2(new_n757), .B1(new_n759), .B2(G1341), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G160), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G29), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n760), .B1(G1341), .B2(new_n759), .C1(new_n761), .C2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n744), .B(new_n768), .C1(new_n741), .C2(new_n743), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n715), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n715), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT29), .Z(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT90), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n694), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT91), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n756), .A2(new_n757), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n767), .A2(new_n761), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n772), .A2(new_n773), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n738), .A2(new_n739), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n694), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n610), .B2(new_n694), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT30), .B(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n715), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n633), .B2(new_n715), .ZN(new_n795));
  NAND2_X1  g370(.A1(G164), .A2(G29), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G27), .B2(G29), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n715), .A2(G33), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT25), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n466), .A2(G139), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n478), .A2(G127), .A3(new_n480), .ZN(new_n806));
  NAND2_X1  g381(.A1(G115), .A2(G2104), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n468), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n801), .B1(new_n809), .B2(new_n715), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2072), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n800), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n715), .A2(G26), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT28), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n487), .A2(G128), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n466), .A2(G140), .ZN(new_n816));
  OR2_X1    g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G29), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT86), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(KEYINPUT86), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2067), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n787), .A2(new_n790), .A3(new_n812), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n734), .A2(new_n769), .A3(new_n782), .A4(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NAND3_X1  g402(.A1(new_n509), .A2(new_n516), .A3(G93), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n516), .A2(G55), .A3(G543), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT93), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT93), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n509), .B2(G67), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n835));
  OAI21_X1  g410(.A(G651), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g411(.A(KEYINPUT92), .B(new_n833), .C1(new_n509), .C2(G67), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n830), .A2(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT94), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n507), .A2(new_n508), .ZN(new_n840));
  INV_X1    g415(.A(new_n504), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n840), .A2(G67), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n832), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT92), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n834), .A2(new_n835), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n845), .A3(G651), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n846), .B(new_n847), .C1(new_n831), .C2(new_n830), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n839), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND3_X1  g426(.A1(new_n839), .A2(new_n613), .A3(new_n848), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n838), .A2(new_n550), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n600), .A2(new_n611), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT38), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n851), .B1(new_n862), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n633), .B(new_n492), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G160), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n819), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n754), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n753), .A2(new_n819), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n501), .A2(new_n500), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT96), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n809), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n809), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n487), .A2(G130), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n466), .A2(G142), .ZN(new_n889));
  OR2_X1    g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n621), .A2(new_n622), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n621), .B2(new_n622), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n893), .A2(new_n894), .A3(new_n721), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n721), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n887), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n887), .A2(KEYINPUT98), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n885), .A2(new_n897), .A3(new_n886), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n868), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n904), .B(KEYINPUT97), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n867), .B(KEYINPUT99), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT40), .B1(new_n907), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G395));
  OAI21_X1  g490(.A(new_n615), .B1(new_n855), .B2(new_n856), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n852), .A2(new_n854), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT95), .ZN(new_n918));
  INV_X1    g493(.A(new_n615), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n600), .A2(G299), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n595), .A2(new_n560), .A3(new_n599), .A4(new_n565), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(KEYINPUT100), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n924), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n928), .A2(KEYINPUT100), .A3(KEYINPUT41), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n916), .A2(new_n921), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n928), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n916), .B2(new_n921), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n916), .A2(new_n921), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n928), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n931), .ZN(new_n939));
  XNOR2_X1  g514(.A(G305), .B(G303), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n591), .ZN(new_n941));
  NAND2_X1  g516(.A1(G290), .A2(G288), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(KEYINPUT101), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n690), .B(G303), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(KEYINPUT101), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n935), .A2(new_n939), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n935), .B2(new_n939), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n849), .A2(new_n605), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n932), .A2(new_n934), .A3(KEYINPUT42), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n938), .B1(new_n937), .B2(new_n931), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n605), .B1(new_n962), .B2(new_n953), .ZN(new_n963));
  INV_X1    g538(.A(new_n958), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT102), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n965), .ZN(G295));
  NAND2_X1  g541(.A1(new_n956), .A2(new_n958), .ZN(G331));
  NOR2_X1   g542(.A1(G168), .A2(G171), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n602), .B2(G168), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n855), .B2(new_n856), .ZN(new_n970));
  INV_X1    g545(.A(new_n968), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(G301), .B2(G286), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n918), .A2(new_n920), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n973), .A3(new_n933), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n970), .A2(new_n973), .A3(KEYINPUT104), .A4(new_n933), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n973), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n925), .A2(KEYINPUT103), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(new_n926), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n952), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n970), .A2(new_n973), .A3(new_n933), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n930), .B1(new_n970), .B2(new_n973), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n986), .B2(new_n951), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n983), .A2(new_n987), .A3(KEYINPUT105), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n974), .A2(new_n975), .B1(new_n978), .B2(new_n980), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n951), .B1(new_n991), .B2(new_n977), .ZN(new_n992));
  INV_X1    g567(.A(new_n930), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n855), .A2(new_n856), .A3(new_n969), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n972), .B1(new_n918), .B2(new_n920), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(new_n951), .A3(new_n974), .ZN(new_n997));
  INV_X1    g572(.A(G37), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n988), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n986), .A2(new_n951), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n989), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT106), .B1(new_n992), .B2(new_n1002), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n983), .A2(new_n987), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1009), .A3(KEYINPUT43), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n999), .A2(new_n1001), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(new_n1013), .ZN(G397));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n877), .A2(new_n1015), .A3(new_n878), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n877), .A2(KEYINPUT107), .A3(new_n1015), .A4(new_n878), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n483), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n467), .A2(new_n473), .B1(G101), .B2(new_n475), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(G40), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n819), .B(G2067), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT109), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n721), .A2(new_n725), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n722), .A2(new_n724), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n753), .B(G1996), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n591), .B(G1986), .Z(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1025), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT112), .B(G8), .Z(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n873), .B2(new_n874), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1019), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G40), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n477), .A2(new_n483), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1043), .B(new_n1045), .C1(KEYINPUT45), .C2(new_n1041), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n742), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1041), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT114), .B(G2084), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1045), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1038), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1037), .B(new_n1040), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT123), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n875), .A2(new_n1015), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1024), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n743), .B1(new_n1062), .B2(new_n1043), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1052), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1047), .A2(new_n1066), .A3(new_n1052), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(G8), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT122), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1065), .A2(new_n1067), .A3(new_n1070), .A4(G8), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1040), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1059), .B1(new_n1072), .B2(KEYINPUT51), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1065), .A2(new_n1039), .A3(new_n1067), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT62), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1071), .A2(new_n1040), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1037), .B1(new_n1078), .B2(new_n1069), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1077), .B(new_n1074), .C1(new_n1079), .C2(new_n1059), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1084), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1086), .A2(KEYINPUT111), .A3(new_n1082), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G8), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n877), .A2(KEYINPUT45), .A3(new_n1015), .A4(new_n878), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1061), .A2(new_n1019), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1045), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n698), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1048), .A2(new_n1050), .A3(new_n1045), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT110), .B(G2090), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1089), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1086), .A2(new_n1082), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1092), .A2(new_n698), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1038), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT49), .ZN(new_n1102));
  OAI21_X1  g677(.A(G1981), .B1(new_n579), .B2(new_n582), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n579), .A2(new_n582), .A3(G1981), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1105), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT49), .A3(new_n1103), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1038), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT113), .B(G1976), .Z(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1112), .B(new_n1109), .C1(new_n1113), .C2(G288), .ZN(new_n1114));
  NAND3_X1  g689(.A1(G160), .A2(G40), .A3(new_n1041), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1054), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(new_n1113), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT52), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1098), .A2(new_n1101), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1090), .A2(new_n798), .A3(new_n1045), .A4(new_n1091), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1048), .A2(new_n1050), .A3(new_n1045), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1122), .A2(new_n1123), .B1(new_n739), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1062), .A2(new_n1043), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n602), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1121), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1076), .A2(new_n1080), .A3(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1110), .A2(new_n1113), .A3(new_n701), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1109), .B1(new_n1133), .B2(new_n1105), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1098), .B2(new_n1119), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1119), .B1(new_n1088), .B2(new_n1097), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1055), .A2(new_n1137), .A3(G286), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1099), .B1(new_n1097), .B2(KEYINPUT115), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1136), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT116), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1055), .A2(G286), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1098), .A2(new_n1143), .A3(new_n1101), .A4(new_n1120), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1141), .A2(new_n1142), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(KEYINPUT116), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1135), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1348), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1115), .B2(G2067), .ZN(new_n1152));
  INV_X1    g727(.A(G2067), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1045), .A2(KEYINPUT118), .A3(new_n1153), .A4(new_n1041), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(new_n610), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n610), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1115), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1996), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1090), .A2(new_n1166), .A3(new_n1045), .A4(new_n1091), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1115), .A2(KEYINPUT120), .A3(new_n1162), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n550), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1172), .A3(new_n550), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1124), .A2(new_n780), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT56), .B(G2072), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1090), .A2(new_n1045), .A3(new_n1091), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT119), .ZN(new_n1181));
  NAND3_X1  g756(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1182));
  OR2_X1    g757(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1183));
  NAND2_X1  g758(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n560), .A2(new_n565), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1180), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n1177), .A3(new_n1175), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1189), .A2(KEYINPUT61), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1189), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1186), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1161), .A2(new_n1174), .A3(new_n1191), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1188), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1155), .A2(new_n610), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1189), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1021), .A2(new_n1045), .A3(new_n1127), .A4(new_n1090), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n567), .B1(new_n1201), .B2(new_n1125), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1125), .A2(G301), .A3(new_n1128), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT54), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1201), .A2(new_n1125), .A3(G301), .ZN(new_n1206));
  AOI21_X1  g781(.A(KEYINPUT54), .B1(new_n1130), .B2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1205), .A2(new_n1207), .A3(new_n1121), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1200), .B(new_n1208), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1148), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1036), .B1(new_n1132), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1025), .B1(new_n753), .B2(new_n1026), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT126), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT47), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1025), .A2(new_n1166), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT46), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1214), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1025), .ZN(new_n1219));
  NOR3_X1   g794(.A1(new_n1219), .A2(G1986), .A3(G290), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT48), .ZN(new_n1221));
  OAI22_X1  g796(.A1(new_n1217), .A2(new_n1218), .B1(new_n1034), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1028), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n869), .A2(new_n1153), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1223), .B1(new_n1226), .B2(new_n1025), .ZN(new_n1227));
  AOI211_X1 g802(.A(KEYINPUT125), .B(new_n1219), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1222), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1211), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g805(.A1(new_n907), .A2(new_n912), .ZN(new_n1232));
  NOR3_X1   g806(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1233));
  AND2_X1   g807(.A1(new_n685), .A2(new_n686), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n685), .A2(new_n686), .ZN(new_n1235));
  OAI21_X1  g809(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1237));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n687), .A2(new_n1238), .A3(new_n1233), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  AND3_X1   g814(.A1(new_n1004), .A2(new_n1232), .A3(new_n1240), .ZN(G308));
  NAND3_X1  g815(.A1(new_n1004), .A2(new_n1232), .A3(new_n1240), .ZN(G225));
endmodule


