//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n209), .B(new_n214), .C1(new_n215), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n215), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT64), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G351));
  NAND3_X1  g0042(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT70), .ZN(new_n244));
  INV_X1    g0044(.A(G77), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT71), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n212), .ZN(new_n249));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(KEYINPUT70), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n249), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n203), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G77), .A3(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT8), .B(G58), .Z(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT15), .B(G87), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n249), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n247), .A2(new_n257), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT72), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n268), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G33), .A3(G41), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(G274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n280), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G244), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G238), .A3(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(G232), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G107), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n289), .B(new_n291), .C1(new_n292), .C2(new_n288), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n276), .A2(new_n272), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n286), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n287), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(G179), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n271), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n269), .A2(new_n270), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n249), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G58), .A2(G68), .ZN(new_n309));
  INV_X1    g0109(.A(G50), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n204), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n311), .B(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n258), .A2(new_n262), .B1(G150), .B2(new_n259), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n308), .A2(new_n243), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n256), .A2(G50), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n316), .A2(new_n317), .B1(G50), .B2(new_n243), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n294), .B1(new_n323), .B2(new_n245), .ZN(new_n324));
  MUX2_X1   g0124(.A(G222), .B(G223), .S(G1698), .Z(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n277), .A2(G226), .A3(new_n282), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n281), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n319), .B1(new_n300), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G179), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n304), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(KEYINPUT9), .B2(new_n319), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT9), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n315), .B2(new_n318), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n336), .A2(KEYINPUT10), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(KEYINPUT10), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n307), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G232), .ZN(new_n341));
  MUX2_X1   g0141(.A(G223), .B(G226), .S(G1698), .Z(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n288), .B1(G33), .B2(G87), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n281), .B1(new_n283), .B2(new_n341), .C1(new_n343), .C2(new_n294), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n304), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G200), .B2(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n258), .A2(new_n256), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n347), .A2(new_n316), .B1(new_n243), .B2(new_n258), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G58), .ZN(new_n350));
  INV_X1    g0150(.A(G68), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n309), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n259), .A2(G159), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT77), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n288), .C2(G20), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT78), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n204), .A2(KEYINPUT7), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n323), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT78), .B1(new_n288), .B2(new_n363), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n323), .A2(new_n204), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n359), .B1(new_n368), .B2(new_n360), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT79), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(G20), .B1(new_n320), .B2(new_n322), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT77), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(new_n361), .A3(new_n366), .A4(new_n365), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT79), .A3(G68), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n358), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n261), .A3(KEYINPUT3), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n364), .C1(new_n323), .C2(new_n378), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n360), .B1(new_n288), .B2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n355), .B1(new_n382), .B2(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n249), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n346), .B(new_n349), .C1(new_n377), .C2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT17), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n375), .A2(KEYINPUT79), .A3(G68), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT79), .B1(new_n375), .B2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n357), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n384), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n348), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n346), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n344), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(G169), .B2(new_n344), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n349), .B1(new_n377), .B2(new_n384), .ZN(new_n401));
  INV_X1    g0201(.A(new_n399), .ZN(new_n402));
  INV_X1    g0202(.A(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n340), .A2(new_n395), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT12), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n244), .B2(new_n351), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT74), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n251), .A2(new_n408), .A3(G20), .A4(new_n351), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n262), .A2(G77), .B1(G20), .B2(new_n351), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n259), .A2(G50), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n308), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XOR2_X1   g0215(.A(new_n415), .B(KEYINPUT11), .Z(new_n416));
  NAND3_X1  g0216(.A1(new_n255), .A2(G68), .A3(new_n256), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n277), .A2(G238), .A3(new_n282), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G226), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n341), .B2(G1698), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n424), .B2(new_n288), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n281), .B(new_n420), .C1(new_n425), .C2(new_n294), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT13), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT73), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n341), .A2(G1698), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G226), .B2(G1698), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n421), .B1(new_n430), .B2(new_n323), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n295), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n281), .A4(new_n420), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n427), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  OR3_X1    g0235(.A1(new_n426), .A2(new_n428), .A3(KEYINPUT13), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(G169), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n438), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(G169), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n427), .A2(G179), .A3(new_n434), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n419), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n443), .ZN(new_n445));
  AOI211_X1 g0245(.A(KEYINPUT76), .B(new_n445), .C1(new_n439), .C2(new_n441), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n418), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n427), .A2(G190), .A3(new_n434), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n412), .A2(new_n448), .A3(new_n416), .A4(new_n417), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n435), .A2(new_n436), .A3(G200), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n407), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n203), .A2(G45), .ZN(new_n454));
  OR2_X1    g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n277), .A3(G274), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n277), .A3(KEYINPUT82), .A4(G274), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n320), .A2(new_n322), .A3(G250), .A4(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n320), .A2(new_n322), .A3(G244), .A4(new_n290), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n295), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n455), .A2(new_n456), .ZN(new_n470));
  INV_X1    g0270(.A(new_n454), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n472), .A2(new_n277), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G257), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n462), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n292), .B1(new_n380), .B2(new_n381), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n259), .A2(G77), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n478), .A2(new_n479), .A3(G107), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n477), .B1(new_n482), .B2(new_n204), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n249), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n243), .A2(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n203), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n243), .A2(new_n486), .A3(new_n212), .A4(new_n248), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(G97), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n475), .A2(new_n300), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n462), .A2(new_n469), .A3(new_n474), .A4(new_n397), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n475), .A2(G200), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n462), .A2(new_n469), .A3(new_n474), .A4(G190), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(new_n484), .A3(new_n489), .A4(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n320), .A2(new_n322), .A3(G257), .A4(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n320), .A2(new_n322), .A3(G250), .A4(new_n290), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n295), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n472), .A2(G264), .A3(new_n277), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT90), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(KEYINPUT90), .A3(new_n502), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(G179), .A3(new_n506), .A4(new_n462), .ZN(new_n507));
  INV_X1    g0307(.A(new_n462), .ZN(new_n508));
  OAI21_X1  g0308(.A(G169), .B1(new_n508), .B2(new_n503), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n320), .A2(new_n322), .A3(new_n204), .A4(G87), .ZN(new_n511));
  AND2_X1   g0311(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n288), .A2(new_n204), .A3(G87), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(G20), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n204), .B2(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n292), .A2(KEYINPUT23), .A3(G20), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT24), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT24), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n515), .A2(new_n516), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n308), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g0327(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n528));
  NOR2_X1   g0328(.A1(new_n243), .A2(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n292), .B2(new_n487), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n510), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n505), .A2(new_n462), .A3(new_n506), .ZN(new_n535));
  INV_X1    g0335(.A(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n508), .A2(new_n503), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n304), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n532), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n496), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n288), .A2(new_n204), .A3(G68), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n262), .A2(G97), .ZN(new_n544));
  AND2_X1   g0344(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n422), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(KEYINPUT84), .A3(new_n204), .ZN(new_n551));
  NOR3_X1   g0351(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT84), .B1(new_n550), .B2(new_n204), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n249), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n244), .A2(new_n264), .ZN(new_n558));
  AOI21_X1  g0358(.A(G250), .B1(new_n203), .B2(G45), .ZN(new_n559));
  INV_X1    g0359(.A(G274), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n471), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n561), .A2(new_n277), .ZN(new_n562));
  OR2_X1    g0362(.A1(G238), .A2(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n284), .A2(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n320), .A2(new_n563), .A3(new_n322), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n294), .B1(new_n565), .B2(new_n517), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n487), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n557), .A2(new_n558), .A3(new_n567), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n558), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n556), .B2(new_n249), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n567), .A4(new_n571), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n565), .A2(new_n517), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n295), .B1(new_n277), .B2(new_n561), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n264), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n488), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n543), .A2(new_n548), .ZN(new_n584));
  XNOR2_X1  g0384(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n585));
  AOI21_X1  g0385(.A(G20), .B1(new_n585), .B2(new_n422), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n552), .B1(new_n586), .B2(KEYINPUT84), .ZN(new_n587));
  INV_X1    g0387(.A(new_n555), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n558), .B(new_n583), .C1(new_n589), .C2(new_n308), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n579), .A2(G169), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n562), .A2(new_n566), .A3(G179), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n581), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(G116), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n203), .B2(G33), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n255), .A2(new_n597), .B1(new_n244), .B2(new_n596), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n463), .B(new_n204), .C1(G33), .C2(new_n479), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n249), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n300), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n473), .A2(G270), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n288), .A2(G257), .A3(new_n290), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n323), .A2(G303), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n295), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n462), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n604), .A2(new_n611), .A3(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n603), .A2(new_n598), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n460), .A2(new_n461), .B1(new_n473), .B2(G270), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(G179), .A4(new_n610), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n611), .B2(G200), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n304), .B2(new_n611), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n604), .A2(new_n611), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT87), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n622), .B(KEYINPUT21), .C1(new_n604), .C2(new_n611), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n616), .B(new_n618), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n542), .A2(new_n595), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n453), .A2(new_n625), .ZN(G372));
  OR2_X1    g0426(.A1(new_n337), .A2(new_n338), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n451), .A2(new_n299), .A3(new_n271), .A4(new_n301), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n394), .B1(new_n447), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT92), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n392), .B2(new_n399), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n401), .A2(KEYINPUT92), .A3(new_n402), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n627), .B1(new_n629), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT93), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(new_n640), .A3(new_n330), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n639), .B2(new_n330), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n453), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n534), .B(new_n616), .C1(new_n621), .C2(new_n623), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n576), .A2(new_n567), .A3(new_n571), .A4(new_n580), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n594), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n532), .B2(new_n540), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n648), .A3(new_n496), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n490), .B2(new_n491), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n647), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n475), .A2(new_n300), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n484), .A2(new_n489), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(new_n491), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n650), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT26), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(KEYINPUT26), .A2(new_n581), .A3(new_n594), .A4(new_n655), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n649), .B(new_n594), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n643), .B1(new_n644), .B2(new_n660), .ZN(G369));
  OAI21_X1  g0461(.A(new_n616), .B1(new_n621), .B2(new_n623), .ZN(new_n662));
  INV_X1    g0462(.A(new_n624), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n251), .A2(new_n204), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT94), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n613), .ZN(new_n671));
  MUX2_X1   g0471(.A(new_n662), .B(new_n663), .S(new_n671), .Z(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n532), .B1(new_n509), .B2(new_n507), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n670), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n532), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n670), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n662), .A2(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n675), .A2(new_n677), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n203), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n553), .A2(G116), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n211), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  NAND2_X1  g0495(.A1(new_n492), .A2(new_n495), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n674), .A2(new_n696), .A3(new_n675), .ZN(new_n697));
  INV_X1    g0497(.A(new_n595), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n663), .A4(new_n677), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n610), .A2(G179), .A3(new_n579), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n614), .A3(new_n505), .A4(new_n506), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT30), .B1(new_n701), .B2(new_n475), .ZN(new_n702));
  AND4_X1   g0502(.A1(G179), .A2(new_n614), .A3(new_n579), .A4(new_n610), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n505), .A2(new_n506), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  INV_X1    g0505(.A(new_n475), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n535), .A2(new_n475), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI211_X1 g0511(.A(G179), .B(new_n579), .C1(new_n614), .C2(new_n610), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n535), .A2(KEYINPUT95), .A3(new_n475), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n677), .B1(new_n715), .B2(KEYINPUT96), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n708), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n699), .A2(KEYINPUT31), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n720), .B(new_n677), .C1(new_n708), .C2(new_n714), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n647), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n492), .A2(KEYINPUT91), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n656), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n726), .A2(KEYINPUT26), .B1(new_n590), .B2(new_n593), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n496), .A2(KEYINPUT97), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT97), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n696), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n728), .A2(new_n645), .A3(new_n648), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n698), .A2(new_n655), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n727), .B(new_n731), .C1(KEYINPUT26), .C2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n660), .A2(new_n670), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n735), .B2(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n695), .B1(new_n738), .B2(G1), .ZN(G364));
  INV_X1    g0539(.A(new_n673), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n250), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT98), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n692), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n672), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n207), .A2(new_n288), .ZN(new_n748));
  INV_X1    g0548(.A(G355), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(G116), .B2(new_n207), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n241), .A2(G45), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n690), .A2(new_n288), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n279), .B2(new_n211), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT99), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n212), .B1(G20), .B2(new_n300), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n745), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n204), .A2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n536), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT102), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G283), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n204), .A2(new_n304), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n397), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G322), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n763), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G329), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n770), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(new_n764), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G303), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n763), .A2(new_n769), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n323), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n204), .B1(new_n772), .B2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(G294), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n204), .A2(new_n397), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n785), .A2(new_n304), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G326), .A2(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n767), .A2(new_n778), .A3(new_n784), .A4(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n766), .A2(G107), .ZN(new_n793));
  INV_X1    g0593(.A(new_n773), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n796));
  OAI221_X1 g0596(.A(new_n288), .B1(new_n568), .B2(new_n776), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n782), .A2(new_n479), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G68), .B2(new_n789), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n770), .ZN(new_n803));
  INV_X1    g0603(.A(new_n779), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G58), .A2(new_n803), .B1(new_n804), .B2(G77), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n310), .B2(new_n786), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n792), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n762), .B1(new_n808), .B2(new_n759), .ZN(new_n809));
  INV_X1    g0609(.A(new_n758), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n672), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n747), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  NOR2_X1   g0613(.A1(new_n307), .A2(new_n670), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n659), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n302), .A2(new_n670), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n271), .A2(new_n670), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n306), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n302), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n815), .B1(new_n735), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n745), .B1(new_n723), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n723), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n759), .A2(new_n756), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n744), .B1(new_n245), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n759), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n288), .B(new_n800), .C1(G107), .C2(new_n777), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n766), .A2(G87), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G283), .A2(new_n789), .B1(new_n787), .B2(G303), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n779), .A2(new_n596), .B1(new_n773), .B2(new_n780), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G294), .B2(new_n803), .ZN(new_n830));
  AND4_X1   g0630(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n788), .A2(new_n832), .B1(new_n786), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT103), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  INV_X1    g0636(.A(G159), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n770), .C1(new_n837), .C2(new_n779), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT104), .Z(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n766), .A2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n288), .B1(new_n773), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G50), .B2(new_n777), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(new_n350), .C2(new_n782), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n839), .B2(KEYINPUT34), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n831), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n824), .B1(new_n819), .B2(new_n757), .C1(new_n825), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n822), .A2(new_n848), .ZN(G384));
  INV_X1    g0649(.A(new_n482), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n850), .A2(KEYINPUT35), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(KEYINPUT35), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(G116), .A3(new_n213), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n854));
  XNOR2_X1  g0654(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n211), .B(G77), .C1(new_n350), .C2(new_n351), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n310), .A2(G68), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n203), .B(G13), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n418), .A2(new_n670), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n447), .A2(new_n451), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n447), .B2(new_n451), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n816), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT106), .B1(new_n815), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT106), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n867), .B(new_n816), .C1(new_n659), .C2(new_n814), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n372), .A2(new_n376), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n308), .B1(new_n871), .B2(new_n357), .ZN(new_n872));
  INV_X1    g0672(.A(new_n355), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n388), .B2(new_n389), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n356), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n348), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n385), .B1(new_n876), .B2(new_n668), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n399), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n668), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n401), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n385), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n392), .B2(new_n399), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n871), .B2(new_n873), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n390), .A2(new_n249), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n349), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n880), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n394), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n886), .A2(KEYINPUT107), .A3(new_n893), .A4(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n882), .A2(new_n884), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(new_n402), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n890), .A2(new_n900), .A3(new_n385), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n901), .B2(KEYINPUT37), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n890), .B1(new_n395), .B2(new_n406), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n870), .A2(new_n905), .B1(new_n638), .B2(new_n668), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT18), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT18), .B1(new_n631), .B2(new_n632), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n395), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n881), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n882), .B1(new_n631), .B2(new_n632), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n885), .B1(new_n912), .B2(new_n883), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n902), .A2(new_n903), .A3(new_n898), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT39), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(KEYINPUT39), .B2(new_n905), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n447), .A2(new_n670), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n906), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n453), .B(new_n734), .C1(new_n735), .C2(KEYINPUT29), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n643), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G330), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n819), .B1(new_n861), .B2(new_n862), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n719), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT40), .B1(new_n905), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n881), .B1(new_n637), .B2(new_n395), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n633), .A2(new_n385), .A3(new_n881), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n899), .B1(new_n931), .B2(KEYINPUT37), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n898), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n929), .B1(new_n933), .B2(new_n894), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n928), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n644), .A2(new_n926), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n923), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n203), .B2(new_n742), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n922), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n859), .B1(new_n940), .B2(new_n941), .ZN(G367));
  OAI21_X1  g0742(.A(new_n760), .B1(new_n207), .B2(new_n264), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n753), .A2(new_n232), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n745), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G50), .A2(new_n804), .B1(new_n794), .B2(G137), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n245), .B2(new_n765), .C1(new_n832), .C2(new_n770), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n288), .B1(new_n776), .B2(new_n350), .C1(new_n837), .C2(new_n788), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n782), .A2(new_n351), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n786), .A2(new_n836), .ZN(new_n950));
  NOR4_X1   g0750(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n804), .A2(G283), .ZN(new_n952));
  INV_X1    g0752(.A(G303), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n952), .B1(new_n479), .B2(new_n765), .C1(new_n953), .C2(new_n770), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n776), .A2(new_n596), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT46), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n786), .A2(new_n780), .B1(new_n782), .B2(new_n292), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  INV_X1    g0758(.A(G294), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n323), .B1(new_n773), .B2(new_n958), .C1(new_n788), .C2(new_n959), .ZN(new_n960));
  NOR4_X1   g0760(.A1(new_n954), .A2(new_n956), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n951), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  AOI21_X1  g0763(.A(new_n945), .B1(new_n963), .B2(new_n759), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n576), .A2(new_n571), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n670), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n724), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n594), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n964), .B1(new_n810), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT108), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n743), .A2(G1), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n696), .B(KEYINPUT97), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n670), .A2(new_n654), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n974), .A2(new_n975), .B1(new_n655), .B2(new_n670), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n687), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n976), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n688), .A2(new_n980), .A3(KEYINPUT45), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n687), .B2(new_n976), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n682), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n683), .A3(new_n984), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n685), .B1(new_n680), .B2(new_n684), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n673), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n738), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n691), .B(KEYINPUT41), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n973), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n976), .A2(new_n685), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n974), .A2(new_n675), .A3(new_n975), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n670), .B1(new_n996), .B2(new_n492), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(KEYINPUT42), .B2(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n969), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT43), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n995), .A2(new_n998), .A3(new_n1001), .A4(new_n1000), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n683), .A2(new_n976), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1006), .B(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n972), .B1(new_n993), .B2(new_n1009), .ZN(G387));
  INV_X1    g0810(.A(KEYINPUT110), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n737), .A2(new_n990), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n990), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n723), .A3(new_n736), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n278), .A3(new_n207), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n229), .A2(new_n279), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT109), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n258), .A2(new_n310), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n693), .B(new_n279), .C1(new_n351), .C2(new_n245), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n752), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1016), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(G107), .B2(new_n207), .C1(new_n693), .C2(new_n748), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n744), .B1(new_n1024), .B2(new_n760), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n776), .A2(new_n245), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n323), .B(new_n1026), .C1(new_n258), .C2(new_n789), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n766), .A2(G97), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n782), .A2(new_n264), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G159), .B2(new_n787), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n770), .A2(new_n310), .B1(new_n773), .B2(new_n832), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G68), .B2(new_n804), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n288), .B1(new_n794), .B2(G326), .ZN(new_n1034));
  INV_X1    g0834(.A(G283), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n776), .A2(new_n959), .B1(new_n782), .B2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G317), .A2(new_n803), .B1(new_n804), .B2(G303), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n780), .B2(new_n788), .C1(new_n771), .C2(new_n786), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n1039), .B2(new_n1038), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1034), .B1(new_n596), .B2(new_n765), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n759), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1025), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n681), .B2(new_n758), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1013), .B2(new_n973), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1011), .B1(new_n1015), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1015), .A2(new_n1011), .A3(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(G393));
  INV_X1    g0853(.A(new_n691), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n987), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n683), .B1(new_n979), .B2(new_n984), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1014), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1054), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n988), .A2(new_n1014), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1057), .A2(new_n973), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n237), .A2(new_n752), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n760), .B1(new_n479), .B2(new_n207), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n745), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n323), .B1(new_n776), .B2(new_n1035), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n779), .A2(new_n959), .B1(new_n773), .B2(new_n771), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n788), .A2(new_n953), .B1(new_n782), .B2(new_n596), .ZN(new_n1068));
  OR4_X1    g0868(.A1(new_n793), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n786), .A2(new_n958), .B1(new_n770), .B2(new_n780), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT52), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n323), .B1(new_n804), .B2(new_n258), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G68), .A2(new_n777), .B1(new_n794), .B2(G143), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n782), .A2(new_n245), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G50), .B2(new_n789), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n827), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n786), .A2(new_n832), .B1(new_n770), .B2(new_n837), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1069), .A2(new_n1071), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1065), .B1(new_n1080), .B2(new_n759), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n980), .B2(new_n810), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1061), .A2(new_n1062), .A3(new_n1082), .ZN(G390));
  NAND3_X1  g0883(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n720), .B1(new_n625), .B2(new_n677), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n716), .A2(new_n718), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n453), .A3(G330), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n920), .B(new_n1088), .C1(new_n641), .C2(new_n642), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n862), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n447), .A2(new_n451), .A3(new_n860), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1092), .A2(new_n1087), .A3(G330), .A4(new_n819), .ZN(new_n1093));
  OAI211_X1 g0893(.A(G330), .B(new_n819), .C1(new_n719), .C2(new_n721), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n863), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n866), .A2(new_n869), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1094), .A2(new_n863), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n818), .A2(new_n302), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n733), .A2(new_n677), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n864), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(G330), .B(new_n819), .C1(new_n719), .C2(new_n925), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n863), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1099), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1089), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1092), .B1(new_n865), .B2(new_n868), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n918), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n905), .A2(KEYINPUT39), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT39), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1102), .A2(new_n1092), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n933), .A2(new_n894), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n918), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1113), .A2(new_n1116), .A3(new_n1099), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1093), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1113), .A2(new_n1116), .A3(new_n1099), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1114), .A2(new_n1115), .A3(new_n918), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n917), .B2(new_n1110), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1120), .B(new_n1107), .C1(new_n1122), .C2(new_n1093), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1119), .A2(new_n691), .A3(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1120), .B(new_n973), .C1(new_n1122), .C2(new_n1093), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n823), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n745), .B1(new_n258), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n288), .B(new_n1074), .C1(G87), .C2(new_n777), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G107), .A2(new_n789), .B1(new_n787), .B2(G283), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n770), .A2(new_n596), .B1(new_n779), .B2(new_n479), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G294), .B2(new_n794), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n841), .A2(new_n1128), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n776), .A2(new_n832), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n288), .B1(new_n770), .B2(new_n842), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G137), .B2(new_n789), .ZN(new_n1136));
  INV_X1    g0936(.A(G125), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n765), .A2(new_n310), .B1(new_n773), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n804), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n787), .A2(G128), .B1(new_n783), .B2(G159), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1134), .A2(new_n1136), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n825), .B1(new_n1132), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1127), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n757), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1124), .A2(new_n1148), .A3(KEYINPUT112), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT112), .B1(new_n1124), .B2(new_n1148), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(G378));
  NAND2_X1  g0951(.A1(new_n905), .A2(new_n927), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n929), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n923), .B1(new_n934), .B2(new_n927), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n668), .A2(new_n319), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n1156));
  NAND2_X1  g0956(.A1(new_n339), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n339), .A2(new_n1156), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1155), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n1157), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1160), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1153), .A2(new_n1154), .A3(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT40), .B1(new_n914), .B2(new_n915), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1092), .A2(new_n1087), .A3(new_n819), .ZN(new_n1173));
  OAI21_X1  g0973(.A(G330), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1171), .B1(new_n1174), .B2(new_n928), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n918), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1146), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1170), .A2(new_n1175), .A3(new_n1177), .A4(new_n906), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1170), .A2(new_n1175), .B1(new_n1177), .B2(new_n906), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n973), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1169), .A2(new_n757), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G33), .A2(G41), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G50), .B(new_n1183), .C1(new_n323), .C2(new_n278), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n803), .A2(G107), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT113), .Z(new_n1186));
  NOR2_X1   g0986(.A1(new_n788), .A2(new_n479), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G116), .B2(new_n787), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n773), .A2(new_n1035), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n765), .A2(new_n350), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n582), .C2(new_n804), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1026), .A2(new_n949), .A3(G41), .A4(new_n288), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1186), .A2(new_n1188), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT58), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1184), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n776), .A2(new_n1139), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT114), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(KEYINPUT114), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G125), .B2(new_n787), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n803), .B1(new_n804), .B2(G137), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n789), .A2(G132), .B1(new_n783), .B2(G150), .ZN(new_n1201));
  AND4_X1   g1001(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1183), .B1(new_n765), .B2(new_n837), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G124), .B2(new_n794), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT59), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1195), .B1(new_n1194), .B2(new_n1193), .C1(new_n1204), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n759), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n745), .C1(G50), .C2(new_n1126), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1182), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1181), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1089), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1123), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1174), .A2(new_n928), .A3(new_n1171), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1169), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n919), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1178), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1219), .B2(new_n1178), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1054), .B1(new_n1224), .B2(new_n1216), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1214), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G375));
  NAND2_X1  g1027(.A1(new_n863), .A2(new_n756), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n745), .B1(G68), .B2(new_n1126), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n776), .A2(new_n479), .B1(new_n773), .B2(new_n953), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT120), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1029), .B(new_n1231), .C1(G283), .C2(new_n803), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n288), .B1(new_n766), .B2(G77), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT119), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n786), .A2(new_n959), .B1(new_n779), .B2(new_n292), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G116), .B2(new_n789), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT118), .Z(new_n1237));
  NAND3_X1  g1037(.A1(new_n1232), .A2(new_n1234), .A3(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT121), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n323), .B(new_n1190), .C1(G50), .C2(new_n783), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G137), .A2(new_n803), .B1(new_n804), .B2(G150), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G159), .A2(new_n777), .B1(new_n794), .B2(G128), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G132), .A2(new_n787), .B1(new_n789), .B2(new_n1140), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1238), .A2(KEYINPUT121), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1239), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1229), .B1(new_n1246), .B2(new_n759), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1228), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1094), .A2(new_n863), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(new_n1102), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1250), .A2(new_n1105), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n973), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1248), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT117), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1254), .A3(new_n1089), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1098), .A2(new_n1089), .A3(new_n1106), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT117), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1108), .A2(new_n992), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1253), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(G381));
  XOR2_X1   g1061(.A(new_n1226), .B(KEYINPUT123), .Z(new_n1262));
  NAND2_X1  g1062(.A1(new_n1124), .A2(new_n1148), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(G381), .A2(G387), .A3(G390), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1051), .A2(new_n812), .A3(new_n1052), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(G384), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1262), .A2(new_n1264), .A3(new_n1265), .A4(new_n1268), .ZN(G407));
  INV_X1    g1069(.A(G213), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(G343), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1262), .A2(new_n1264), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G407), .A2(G213), .A3(new_n1272), .ZN(G409));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1266), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1062), .A2(new_n1082), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G387), .A2(KEYINPUT125), .A3(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G390), .B(new_n972), .C1(new_n993), .C2(new_n1009), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT125), .B1(G387), .B2(new_n1278), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1276), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G387), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1284), .B2(G390), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G387), .A2(new_n1286), .A3(new_n1278), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1285), .A2(new_n1275), .A3(new_n1280), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(G384), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n691), .B1(new_n1256), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1258), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1291), .B1(new_n1295), .B2(new_n1253), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1255), .B(new_n1257), .C1(new_n1292), .C2(new_n1107), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1293), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1253), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(G384), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1271), .A2(G2897), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1296), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1302), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1291), .B(new_n1253), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1216), .A2(new_n1220), .A3(new_n992), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n973), .B1(new_n1220), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT124), .B1(new_n1219), .B2(new_n1178), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1213), .B(new_n1309), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(G378), .A2(new_n1226), .B1(new_n1264), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1308), .B1(new_n1314), .B2(new_n1271), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1216), .A2(new_n1220), .A3(KEYINPUT57), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1215), .A2(new_n1123), .B1(new_n1219), .B2(new_n1178), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1318), .B(new_n691), .C1(KEYINPUT57), .C2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT112), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1263), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1124), .A2(new_n1148), .A3(KEYINPUT112), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1214), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(new_n1322), .A3(new_n1323), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1313), .A2(new_n1264), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1271), .B(new_n1317), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1315), .B(new_n1316), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1271), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1296), .A4(new_n1301), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1332), .A2(KEYINPUT62), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1290), .B1(new_n1329), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1290), .B1(new_n1332), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1327), .A2(KEYINPUT63), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1336), .A2(new_n1316), .A3(new_n1337), .A4(new_n1315), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1338), .ZN(G405));
  XNOR2_X1  g1139(.A(new_n1289), .B(new_n1317), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(G375), .A2(new_n1341), .A3(new_n1264), .ZN(new_n1342));
  OAI21_X1  g1142(.A(KEYINPUT127), .B1(new_n1226), .B2(new_n1263), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(new_n1325), .A3(new_n1343), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1340), .B(new_n1344), .ZN(G402));
endmodule


