//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1107, new_n1108;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g021(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n471), .B2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(G2104), .ZN(new_n481));
  OAI211_X1 g056(.A(G137), .B(new_n478), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G101), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n467), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n477), .A2(new_n485), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n470), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n490), .A2(new_n478), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(G136), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(G124), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT69), .ZN(G162));
  NAND4_X1  g073(.A1(new_n490), .A2(G138), .A3(new_n467), .A4(new_n478), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(new_n467), .A3(KEYINPUT71), .A4(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(KEYINPUT71), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(new_n465), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n490), .A2(G126), .A3(G2105), .A4(new_n478), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(new_n467), .B2(G114), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n510));
  OR2_X1    g085(.A1(G102), .A2(G2105), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(G2104), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n525), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AOI22_X1  g105(.A1(new_n519), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n523), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(new_n520), .B1(new_n533), .B2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  XNOR2_X1  g113(.A(KEYINPUT72), .B(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n540), .B1(new_n521), .B2(new_n541), .C1(new_n542), .C2(new_n527), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(G171));
  XOR2_X1   g119(.A(KEYINPUT73), .B(G81), .Z(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n521), .A2(new_n545), .B1(new_n523), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n533), .A2(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(new_n521), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G91), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n559), .B(new_n561), .C1(new_n527), .C2(new_n562), .ZN(G299));
  XNOR2_X1  g138(.A(new_n543), .B(KEYINPUT75), .ZN(G301));
  NAND2_X1  g139(.A1(new_n560), .A2(G87), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n533), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  AOI22_X1  g143(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n527), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n520), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n519), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n527), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT76), .Z(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n560), .A2(G85), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n533), .A2(G47), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n519), .A2(G92), .A3(new_n520), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  AOI22_X1  g161(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n527), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n533), .A2(G54), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n584), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n584), .B1(new_n591), .B2(G868), .ZN(G321));
  MUX2_X1   g168(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g169(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n591), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n591), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n496), .A2(G123), .ZN(new_n602));
  INV_X1    g177(.A(new_n492), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G135), .ZN(new_n604));
  NOR2_X1   g179(.A1(G99), .A2(G2105), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n602), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(G2096), .Z(new_n608));
  NAND3_X1  g183(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(G2100), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(G156));
  XNOR2_X1  g188(.A(G2451), .B(G2454), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT16), .ZN(new_n615));
  XOR2_X1   g190(.A(G2443), .B(G2446), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G1341), .B(G1348), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT77), .B(G2438), .Z(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n619), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G14), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT78), .Z(G401));
  XOR2_X1   g203(.A(G2084), .B(G2090), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2072), .B(G2078), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT79), .ZN(new_n632));
  XOR2_X1   g207(.A(G2067), .B(G2678), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n632), .B(KEYINPUT17), .Z(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n632), .A2(new_n634), .A3(new_n629), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT18), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(new_n633), .A3(new_n629), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2096), .B(G2100), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(G227));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  XOR2_X1   g223(.A(G1956), .B(G2474), .Z(new_n649));
  XOR2_X1   g224(.A(G1961), .B(G1966), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n653));
  INV_X1    g228(.A(new_n648), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n652), .A2(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n648), .A3(new_n651), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n656), .B(new_n658), .C1(new_n652), .C2(new_n653), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1986), .B(G1996), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G1981), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G1991), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G229));
  INV_X1    g240(.A(G29), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G25), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n496), .A2(G119), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  OR2_X1    g244(.A1(G95), .A2(G2105), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n670), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n603), .A2(G131), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n667), .B1(new_n674), .B2(new_n666), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT35), .B(G1991), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  AND2_X1   g254(.A1(KEYINPUT85), .A2(G16), .ZN(new_n680));
  NOR2_X1   g255(.A1(KEYINPUT85), .A2(G16), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n582), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G24), .B2(new_n683), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n677), .B(new_n678), .C1(new_n679), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n683), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G6), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n574), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT86), .Z(new_n694));
  AOI21_X1  g269(.A(new_n689), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(KEYINPUT87), .B1(G16), .B2(G23), .ZN(new_n696));
  OR3_X1    g271(.A1(KEYINPUT87), .A2(G16), .A3(G23), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n696), .B(new_n697), .C1(G288), .C2(new_n691), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n695), .B(new_n700), .C1(new_n690), .C2(new_n694), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT88), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n686), .B1(new_n702), .B2(KEYINPUT34), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n685), .A2(new_n679), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n703), .B(new_n704), .C1(KEYINPUT34), .C2(new_n702), .ZN(new_n705));
  NOR2_X1   g280(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n666), .A2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n603), .A2(G141), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n496), .A2(G129), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT26), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n709), .A2(new_n710), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n708), .B1(new_n715), .B2(new_n666), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT27), .B(G1996), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n705), .A2(new_n706), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n666), .A2(G27), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G164), .B2(new_n666), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2078), .ZN(new_n723));
  NAND2_X1  g298(.A1(G299), .A2(G16), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n683), .A2(KEYINPUT23), .A3(G20), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n726));
  INV_X1    g301(.A(G20), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n682), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1956), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT24), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G34), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(new_n734), .B(G160), .S(G29), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n723), .B(new_n730), .C1(G2084), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n691), .A2(G4), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n591), .B2(new_n691), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT90), .B(G1348), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n607), .A2(new_n666), .ZN(new_n742));
  NAND2_X1  g317(.A1(G171), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G5), .B2(G16), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n746), .B1(new_n745), .B2(new_n744), .C1(new_n736), .C2(G2084), .ZN(new_n747));
  NAND2_X1  g322(.A1(G168), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G21), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n683), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n550), .B2(new_n683), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1341), .Z(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT30), .B2(new_n756), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n751), .A2(new_n752), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n741), .A2(new_n747), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n749), .A2(new_n750), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT25), .Z(new_n763));
  AOI22_X1  g338(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  INV_X1    g339(.A(G139), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n763), .B1(new_n467), .B2(new_n764), .C1(new_n492), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT93), .ZN(new_n767));
  MUX2_X1   g342(.A(G33), .B(new_n767), .S(G29), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2072), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n737), .A2(new_n760), .A3(new_n761), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G35), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G162), .B2(G29), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT29), .Z(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n666), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n496), .A2(G128), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n603), .A2(G140), .ZN(new_n780));
  NOR2_X1   g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n787), .A2(KEYINPUT92), .A3(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT92), .B1(new_n787), .B2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n778), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n770), .A2(new_n775), .A3(new_n776), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n707), .A2(new_n719), .A3(new_n720), .A4(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(G311));
  XNOR2_X1  g369(.A(new_n793), .B(KEYINPUT95), .ZN(G150));
  XOR2_X1   g370(.A(KEYINPUT97), .B(G860), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT96), .B(G93), .Z(new_n797));
  INV_X1    g372(.A(G55), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n521), .A2(new_n797), .B1(new_n523), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n527), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n796), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT37), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n591), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n799), .A2(new_n801), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n550), .B(new_n806), .Z(new_n807));
  XOR2_X1   g382(.A(new_n805), .B(new_n807), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT39), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n796), .B1(new_n810), .B2(KEYINPUT98), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(KEYINPUT98), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(KEYINPUT39), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n803), .B1(new_n812), .B2(new_n813), .ZN(G145));
  XNOR2_X1  g389(.A(G162), .B(new_n607), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G160), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n610), .ZN(new_n817));
  INV_X1    g392(.A(G142), .ZN(new_n818));
  NOR2_X1   g393(.A1(G106), .A2(G2105), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n492), .A2(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G130), .B2(new_n496), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n817), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n787), .B(new_n673), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n714), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n767), .A2(KEYINPUT100), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n505), .A2(new_n827), .A3(new_n514), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n499), .A2(KEYINPUT4), .B1(new_n465), .B2(new_n503), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT99), .B1(new_n829), .B2(new_n513), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n825), .B(new_n832), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n823), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n591), .B1(new_n838), .B2(G299), .ZN(new_n839));
  AND2_X1   g414(.A1(G299), .A2(new_n838), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n598), .B(new_n807), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n841), .B(KEYINPUT41), .Z(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(new_n843), .ZN(new_n846));
  XNOR2_X1  g421(.A(G303), .B(G288), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G305), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n582), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT42), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n846), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G868), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G868), .B2(new_n806), .ZN(G295));
  OAI21_X1  g428(.A(new_n852), .B1(G868), .B2(new_n806), .ZN(G331));
  NOR2_X1   g429(.A1(G168), .A2(new_n543), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G301), .B2(G168), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n807), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n842), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n845), .B2(new_n857), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(new_n849), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n849), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n835), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT43), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n860), .A2(new_n864), .A3(new_n835), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(KEYINPUT102), .ZN(new_n868));
  MUX2_X1   g443(.A(new_n866), .B(new_n868), .S(KEYINPUT44), .Z(G397));
  INV_X1    g444(.A(G1384), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n831), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT45), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n831), .A2(new_n874), .A3(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT67), .B1(new_n475), .B2(G2105), .ZN(new_n877));
  AOI211_X1 g452(.A(new_n464), .B(new_n467), .C1(new_n473), .C2(new_n474), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n485), .B(G40), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G2067), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n787), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n882), .B2(new_n715), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT127), .Z(new_n884));
  NOR2_X1   g459(.A1(new_n880), .A2(G1996), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT46), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT47), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n673), .B(new_n676), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT105), .Z(new_n890));
  INV_X1    g465(.A(G1996), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n714), .B(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n880), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n880), .A2(G1986), .A3(G290), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT48), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n676), .A3(new_n674), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n785), .A2(new_n881), .A3(new_n786), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n880), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n888), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  AOI211_X1 g476(.A(new_n873), .B(G1384), .C1(new_n828), .C2(new_n830), .ZN(new_n902));
  INV_X1    g477(.A(new_n879), .ZN(new_n903));
  AOI21_X1  g478(.A(G1384), .B1(new_n505), .B2(new_n514), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(KEYINPUT45), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT106), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G2078), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n827), .B1(new_n505), .B2(new_n514), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n829), .A2(KEYINPUT99), .A3(new_n513), .ZN(new_n909));
  OAI211_X1 g484(.A(KEYINPUT45), .B(new_n870), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n870), .B1(new_n829), .B2(new_n513), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n879), .B1(new_n873), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n907), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT53), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT50), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n879), .B1(new_n904), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT50), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n912), .B2(KEYINPUT50), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g501(.A(KEYINPUT114), .B(new_n920), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT119), .B(G1961), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n913), .B1(new_n873), .B2(new_n912), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n930), .A2(new_n916), .A3(G2078), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT120), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n918), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT121), .B1(new_n936), .B2(G301), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n929), .A2(new_n934), .A3(new_n931), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n934), .B1(new_n929), .B2(new_n931), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n917), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT121), .ZN(new_n941));
  INV_X1    g516(.A(G301), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n930), .A2(new_n750), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT111), .B(G2084), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n924), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(G8), .ZN(new_n949));
  NAND2_X1  g524(.A1(G286), .A2(G8), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT51), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(G8), .C1(new_n948), .C2(G286), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT118), .ZN(new_n954));
  INV_X1    g529(.A(new_n950), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n948), .A2(new_n954), .A3(new_n955), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n951), .B(new_n953), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(G8), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT55), .Z(new_n963));
  OAI21_X1  g538(.A(KEYINPUT108), .B1(new_n924), .B2(G2090), .ZN(new_n964));
  INV_X1    g539(.A(new_n923), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT50), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n774), .A4(new_n920), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1971), .B1(new_n906), .B2(new_n914), .ZN(new_n971));
  OAI211_X1 g546(.A(G8), .B(new_n963), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n879), .A2(new_n912), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G288), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G1976), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(G8), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT52), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n979));
  INV_X1    g554(.A(G1981), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n574), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n574), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n983), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(KEYINPUT49), .A3(new_n981), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n984), .A2(new_n986), .A3(G8), .A4(new_n974), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n974), .A2(new_n976), .A3(G8), .A4(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n978), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n972), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n920), .B1(new_n919), .B2(new_n904), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(G2090), .ZN(new_n994));
  OAI21_X1  g569(.A(G8), .B1(new_n971), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n963), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n944), .A2(new_n961), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n944), .A2(KEYINPUT125), .A3(new_n961), .A4(new_n998), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1001), .B(new_n1002), .C1(new_n960), .C2(new_n959), .ZN(new_n1003));
  OAI211_X1 g578(.A(G301), .B(new_n917), .C1(new_n938), .C2(new_n939), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n902), .A2(new_n916), .A3(G2078), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n475), .B2(G2105), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n876), .A2(new_n1005), .A3(new_n485), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n917), .A2(new_n929), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G171), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(KEYINPUT54), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT123), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT123), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1004), .A2(new_n1013), .A3(KEYINPUT54), .A4(new_n1010), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n917), .A2(G301), .A3(new_n929), .A4(new_n1008), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT122), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n937), .A2(new_n1018), .A3(new_n943), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n958), .A2(new_n997), .A3(new_n992), .ZN(new_n1022));
  NAND2_X1  g597(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT116), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n550), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT58), .B(G1341), .Z(new_n1027));
  NOR2_X1   g602(.A1(new_n973), .A2(KEYINPUT113), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n903), .A2(KEYINPUT113), .A3(new_n904), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n910), .A2(new_n891), .A3(new_n913), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1026), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1025), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(G299), .B(KEYINPUT57), .Z(new_n1035));
  NOR2_X1   g610(.A1(new_n902), .A2(new_n905), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  INV_X1    g612(.A(G1956), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1036), .A2(new_n1037), .B1(new_n1038), .B2(new_n993), .ZN(new_n1039));
  NAND2_X1  g614(.A1(KEYINPUT117), .A2(KEYINPUT61), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1032), .A2(new_n1033), .A3(new_n1025), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT117), .A3(KEYINPUT61), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n881), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n926), .A2(new_n927), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(G1348), .ZN(new_n1050));
  INV_X1    g625(.A(new_n591), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n591), .B(new_n1048), .C1(new_n1049), .C2(G1348), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(KEYINPUT60), .A3(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1053), .A2(KEYINPUT60), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1044), .A2(new_n1046), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1050), .A2(new_n591), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1045), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1022), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1015), .A2(new_n1021), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n948), .A2(G8), .A3(G168), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n970), .B2(new_n971), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1063), .B(new_n1064), .C1(new_n1065), .C2(new_n996), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1064), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n997), .A2(new_n972), .A3(new_n1067), .A4(new_n991), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n992), .A2(new_n1066), .B1(new_n1068), .B2(new_n1063), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n911), .B1(new_n910), .B2(new_n913), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(new_n964), .A3(new_n969), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1074), .A2(G8), .A3(new_n963), .A4(new_n991), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n984), .A2(new_n986), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n975), .A2(new_n988), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT109), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n981), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(G8), .A3(new_n974), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1075), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1076), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1062), .B1(new_n1069), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1068), .A2(new_n1063), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1063), .B1(new_n1065), .B2(new_n996), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n992), .A2(new_n1067), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1083), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1075), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1092), .A3(KEYINPUT112), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1061), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1061), .B2(new_n1094), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1003), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n880), .A2(new_n679), .A3(new_n582), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n895), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT104), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n894), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1098), .A2(KEYINPUT126), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT126), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n901), .B1(new_n1103), .B2(new_n1104), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g680(.A1(G229), .A2(new_n462), .ZN(new_n1107));
  NOR2_X1   g681(.A1(G401), .A2(G227), .ZN(new_n1108));
  NAND4_X1  g682(.A1(new_n836), .A2(new_n866), .A3(new_n1107), .A4(new_n1108), .ZN(G225));
  INV_X1    g683(.A(G225), .ZN(G308));
endmodule


