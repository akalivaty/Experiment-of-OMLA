//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n217), .A2(new_n227), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  OR2_X1    g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  AOI21_X1  g0047(.A(G1698), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G222), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n249), .B1(new_n250), .B2(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n256), .A3(G274), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(new_n259), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n256), .A2(new_n264), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n258), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n213), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n274), .A2(new_n275), .B1(new_n202), .B2(new_n271), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n207), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(G20), .B2(new_n203), .ZN(new_n283));
  INV_X1    g0083(.A(new_n273), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n268), .A2(G200), .B1(new_n269), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(KEYINPUT9), .B(new_n276), .C1(new_n283), .C2(new_n284), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT67), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n268), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT10), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n268), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n258), .A2(new_n294), .A3(new_n267), .A4(new_n261), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n285), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT66), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n248), .A2(G232), .ZN(new_n299));
  INV_X1    g0099(.A(G107), .ZN(new_n300));
  INV_X1    g0100(.A(G238), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n299), .B1(new_n300), .B2(new_n251), .C1(new_n301), .C2(new_n252), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n257), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n266), .A2(G244), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n261), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(G179), .ZN(new_n306));
  INV_X1    g0106(.A(new_n277), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n284), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n206), .A2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n274), .A2(G77), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G77), .B2(new_n270), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n305), .B2(new_n292), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n314), .A2(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n305), .B2(G200), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n303), .A2(G190), .A3(new_n261), .A4(new_n304), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n306), .A2(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n291), .A2(new_n298), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n281), .A2(new_n202), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n278), .A2(new_n250), .B1(new_n207), .B2(G68), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n273), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT11), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT71), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT72), .B1(new_n271), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT12), .Z(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n206), .B2(G20), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n274), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n330), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n231), .A2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n251), .B(new_n340), .C1(G226), .C2(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT68), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(G33), .A3(G97), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n256), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n301), .B1(new_n263), .B2(new_n265), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  INV_X1    g0150(.A(new_n261), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n256), .A2(new_n264), .A3(new_n259), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n264), .B1(new_n256), .B2(new_n259), .ZN(new_n354));
  OAI21_X1  g0154(.A(G238), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT69), .B1(new_n355), .B2(new_n261), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n339), .B(new_n348), .C1(new_n352), .C2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n348), .B1(new_n352), .B2(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT13), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(KEYINPUT69), .A3(new_n261), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT70), .A3(new_n339), .A4(new_n348), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n359), .A2(new_n361), .A3(G179), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n366), .B(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n292), .B1(new_n361), .B2(new_n357), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT14), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n338), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT77), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G58), .B2(G68), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n246), .A2(new_n207), .A3(new_n247), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n246), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n247), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n376), .B1(new_n381), .B2(G68), .ZN(new_n382));
  AOI211_X1 g0182(.A(KEYINPUT76), .B(new_n332), .C1(new_n379), .C2(new_n380), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT16), .B(new_n375), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n372), .B(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n201), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n207), .B1(new_n389), .B2(new_n281), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n332), .B1(new_n379), .B2(new_n380), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n384), .A2(new_n392), .A3(new_n273), .ZN(new_n393));
  INV_X1    g0193(.A(new_n274), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n307), .A2(new_n315), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n394), .A2(new_n395), .B1(new_n270), .B2(new_n307), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n253), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n251), .B(new_n400), .C1(G226), .C2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n256), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n261), .B1(new_n231), .B2(new_n262), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n292), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n403), .A2(new_n404), .A3(new_n294), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n405), .A2(new_n289), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(G200), .B2(new_n405), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n393), .A2(new_n397), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n408), .B1(new_n393), .B2(new_n397), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n393), .A2(new_n397), .A3(new_n413), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n411), .A2(new_n415), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  OR3_X1    g0222(.A1(new_n324), .A2(new_n371), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n359), .A2(new_n361), .A3(G190), .A4(new_n365), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n339), .B1(new_n364), .B2(new_n348), .ZN(new_n425));
  AOI211_X1 g0225(.A(KEYINPUT13), .B(new_n347), .C1(new_n362), .C2(new_n363), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n338), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT73), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n361), .A2(new_n357), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n337), .B1(new_n430), .B2(G200), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n424), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(KEYINPUT74), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT74), .B1(new_n429), .B2(new_n433), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n423), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(KEYINPUT3), .A2(G33), .ZN(new_n439));
  NOR2_X1   g0239(.A1(KEYINPUT3), .A2(G33), .ZN(new_n440));
  OAI211_X1 g0240(.A(G257), .B(G1698), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(G250), .B(new_n399), .C1(new_n439), .C2(new_n440), .ZN(new_n442));
  INV_X1    g0242(.A(G294), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n311), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n257), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n206), .A2(G45), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  INV_X1    g0247(.A(G41), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT5), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n257), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G264), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n450), .B1(KEYINPUT78), .B2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n256), .A2(G274), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n256), .A2(G274), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT79), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n292), .B1(new_n455), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n257), .A2(new_n444), .B1(new_n453), .B2(G264), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n461), .A3(new_n456), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT79), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n294), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT81), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n475), .B(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n207), .B(G87), .C1(new_n439), .C2(new_n440), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n475), .B(KEYINPUT82), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT23), .B1(new_n300), .B2(G20), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n300), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n484), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n484), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n273), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT25), .B1(new_n271), .B2(new_n300), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n271), .A2(KEYINPUT25), .A3(new_n300), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n311), .A2(G1), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n271), .A2(new_n273), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n496), .A2(new_n497), .B1(new_n499), .B2(G107), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n473), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n471), .A2(new_n445), .A3(new_n454), .A4(new_n289), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT83), .ZN(new_n504));
  INV_X1    g0304(.A(G200), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n455), .B2(new_n466), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n503), .A2(KEYINPUT83), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n494), .B(new_n500), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G264), .B(G1698), .C1(new_n439), .C2(new_n440), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n251), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n439), .A2(new_n440), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G303), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n251), .A2(G257), .A3(new_n399), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n294), .B1(new_n518), .B2(new_n257), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n469), .A2(new_n470), .B1(new_n453), .B2(G270), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n207), .C1(G33), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G20), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n273), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n273), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n270), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n499), .B2(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n519), .A2(new_n520), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n518), .A2(new_n257), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n520), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n292), .B1(new_n530), .B2(new_n532), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n537), .A2(new_n289), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n505), .B1(new_n520), .B2(new_n536), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n543), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n256), .A2(G274), .A3(new_n459), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n256), .A2(G250), .A3(new_n446), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(G1698), .C1(new_n439), .C2(new_n440), .ZN(new_n550));
  OAI211_X1 g0350(.A(G238), .B(new_n399), .C1(new_n439), .C2(new_n440), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n486), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n257), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G169), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n257), .ZN(new_n555));
  INV_X1    g0355(.A(new_n549), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n555), .A2(new_n294), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n310), .A2(new_n270), .ZN(new_n559));
  INV_X1    g0359(.A(G87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n522), .A3(new_n300), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n343), .B2(new_n345), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n563), .B2(G20), .ZN(new_n564));
  AOI21_X1  g0364(.A(G20), .B1(new_n246), .B2(new_n247), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n312), .A2(G97), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n565), .A2(G68), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n559), .B1(new_n568), .B2(new_n273), .ZN(new_n569));
  INV_X1    g0369(.A(new_n499), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n309), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n270), .A2(G97), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n499), .B2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n300), .B1(new_n379), .B2(new_n380), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g0377(.A(G97), .B(G107), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT6), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n579), .A2(new_n522), .A3(G107), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n575), .B1(new_n585), .B2(new_n273), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n469), .A2(new_n470), .B1(new_n453), .B2(G257), .ZN(new_n587));
  OAI211_X1 g0387(.A(G250), .B(G1698), .C1(new_n439), .C2(new_n440), .ZN(new_n588));
  OAI211_X1 g0388(.A(G244), .B(new_n399), .C1(new_n439), .C2(new_n440), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n521), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT4), .B1(new_n248), .B2(G244), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n257), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n586), .B(new_n595), .C1(new_n289), .C2(new_n594), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n581), .B1(new_n579), .B2(new_n578), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n597), .A2(new_n207), .B1(new_n250), .B2(new_n281), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n273), .B1(new_n598), .B2(new_n576), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n594), .A2(new_n292), .B1(new_n599), .B2(new_n574), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n587), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n294), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n555), .A2(new_n556), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n499), .A2(G87), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n555), .A2(G190), .A3(new_n556), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n569), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n572), .A2(new_n596), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n438), .A2(new_n510), .A3(new_n546), .A4(new_n609), .ZN(G372));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n604), .A2(KEYINPUT84), .A3(G200), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n553), .B2(new_n505), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n569), .A2(new_n606), .A3(new_n607), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n571), .B2(new_n558), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n509), .A2(new_n617), .A3(new_n603), .A4(new_n596), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n535), .B(new_n621), .C1(new_n540), .C2(new_n541), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n501), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n619), .B1(new_n623), .B2(KEYINPUT86), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n518), .A2(new_n257), .ZN(new_n625));
  INV_X1    g0425(.A(G270), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n463), .A2(new_n256), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n462), .A2(new_n465), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n539), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n621), .B1(new_n632), .B2(new_n535), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT85), .B(new_n534), .C1(new_n630), .C2(new_n631), .ZN(new_n634));
  OAI211_X1 g0434(.A(KEYINPUT86), .B(new_n502), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n611), .B1(new_n624), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n572), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n572), .A2(new_n600), .A3(new_n608), .A4(new_n602), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n594), .A2(G179), .ZN(new_n642));
  AOI21_X1  g0442(.A(G169), .B1(new_n587), .B2(new_n593), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n642), .A2(new_n586), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n617), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT88), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n640), .A2(KEYINPUT88), .A3(new_n645), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n502), .B1(new_n633), .B2(new_n634), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(KEYINPUT87), .A3(new_n635), .A4(new_n619), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n637), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n438), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n415), .A2(new_n421), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n306), .A2(new_n319), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n429), .B2(new_n433), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n371), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n411), .A2(new_n418), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n297), .B1(new_n661), .B2(new_n291), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(G369));
  NAND3_X1  g0463(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n533), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n546), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n620), .A2(new_n622), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n670), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT89), .Z(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n510), .ZN(new_n676));
  INV_X1    g0476(.A(new_n669), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n494), .B2(new_n500), .ZN(new_n678));
  OAI22_X1  g0478(.A1(new_n676), .A2(new_n678), .B1(new_n502), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n632), .B2(new_n535), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n510), .A2(new_n681), .B1(new_n501), .B2(new_n677), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n210), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n561), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n215), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g0489(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n690));
  XNOR2_X1  g0490(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n501), .A2(new_n542), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n618), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n572), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n641), .B1(new_n617), .B2(new_n644), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n568), .A2(new_n273), .ZN(new_n698));
  INV_X1    g0498(.A(new_n559), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n698), .A2(new_n699), .A3(new_n606), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n607), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n612), .A2(new_n614), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n572), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT26), .B1(new_n703), .B2(new_n603), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n644), .A2(new_n641), .A3(new_n572), .A4(new_n608), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(KEYINPUT92), .A3(new_n572), .A4(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n693), .B1(new_n697), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n669), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n648), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n646), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n624), .A2(new_n636), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(KEYINPUT87), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n669), .B1(new_n715), .B2(new_n637), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n711), .B1(new_n716), .B2(KEYINPUT29), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT91), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n601), .A2(new_n519), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n468), .A2(new_n520), .A3(new_n553), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n718), .B(new_n723), .C1(new_n719), .C2(new_n720), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n601), .B1(new_n471), .B2(new_n468), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n294), .A3(new_n537), .A4(new_n604), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n669), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n510), .A2(new_n609), .A3(new_n546), .A4(new_n677), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n717), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n691), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n206), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n685), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n675), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n674), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n213), .B1(G20), .B2(new_n292), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n207), .B1(new_n747), .B2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n522), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n207), .A2(new_n289), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n505), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G58), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(G179), .A3(new_n505), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n251), .B1(new_n752), .B2(new_n560), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G190), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n749), .B(new_n755), .C1(G68), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(G190), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT96), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(new_n761), .A3(new_n747), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n389), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n756), .A2(new_n289), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT95), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n756), .A2(KEYINPUT95), .A3(new_n289), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G50), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n760), .A2(new_n761), .A3(new_n751), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n300), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n759), .A2(G179), .A3(new_n505), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n773), .B1(new_n779), .B2(G77), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n758), .A2(new_n764), .A3(new_n771), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n772), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n779), .A2(G311), .B1(new_n782), .B2(G283), .ZN(new_n783));
  INV_X1    g0583(.A(new_n762), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G329), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n770), .A2(G326), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n515), .B1(new_n754), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n757), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(new_n443), .B2(new_n748), .ZN(new_n791));
  INV_X1    g0591(.A(new_n752), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n788), .B(new_n791), .C1(G303), .C2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n783), .A2(new_n785), .A3(new_n786), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n746), .B1(new_n781), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n742), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n684), .A2(new_n251), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n244), .A2(new_n458), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n458), .C2(new_n216), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n210), .A2(new_n251), .ZN(new_n801));
  INV_X1    g0601(.A(G355), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n802), .B1(G116), .B2(new_n210), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n800), .B1(KEYINPUT93), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(KEYINPUT93), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n745), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n795), .B(new_n796), .C1(new_n805), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n808), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n673), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n744), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  INV_X1    g0614(.A(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n320), .A2(new_n669), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n323), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n323), .B2(new_n816), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n677), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n653), .A2(new_n649), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n618), .B1(new_n650), .B2(new_n651), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT87), .B1(new_n822), .B2(new_n635), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n817), .A2(new_n818), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n306), .A2(new_n319), .A3(new_n669), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n716), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n742), .B1(new_n828), .B2(new_n735), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n735), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n745), .A2(new_n806), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n742), .B1(G77), .B2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT97), .Z(new_n834));
  OAI221_X1 g0634(.A(new_n251), .B1(new_n748), .B2(new_n753), .C1(new_n202), .C2(new_n752), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G68), .B2(new_n782), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  INV_X1    g0637(.A(G143), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n279), .A2(new_n789), .B1(new_n754), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n769), .A2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(new_n779), .C2(G159), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n836), .B1(new_n837), .B2(new_n762), .C1(new_n842), .C2(KEYINPUT34), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n842), .A2(KEYINPUT34), .ZN(new_n844));
  INV_X1    g0644(.A(G311), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n560), .A2(new_n772), .B1(new_n762), .B2(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n515), .B1(new_n752), .B2(new_n300), .C1(new_n443), .C2(new_n754), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n846), .A2(new_n749), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n769), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n778), .A2(new_n524), .B1(new_n851), .B2(new_n789), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT98), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n843), .A2(new_n844), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT99), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n745), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(KEYINPUT99), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n834), .B1(new_n856), .B2(new_n857), .C1(new_n827), .C2(new_n807), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n830), .A2(new_n858), .ZN(G384));
  NAND2_X1  g0659(.A1(new_n214), .A2(G116), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n583), .B2(KEYINPUT35), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(KEYINPUT35), .B2(new_n583), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT36), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n387), .A2(new_n250), .A3(new_n215), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(G50), .B2(new_n332), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n867));
  OAI211_X1 g0667(.A(G1), .B(new_n738), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT102), .Z(new_n870));
  NOR2_X1   g0670(.A1(new_n657), .A2(new_n669), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n654), .B2(new_n820), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n368), .A2(new_n370), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n337), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n338), .A2(new_n677), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n429), .B2(new_n433), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT74), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n432), .B1(new_n431), .B2(new_n424), .ZN(new_n879));
  AND4_X1   g0679(.A1(new_n432), .A2(new_n424), .A3(new_n338), .A4(new_n427), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n873), .B1(new_n881), .B2(new_n434), .ZN(new_n882));
  INV_X1    g0682(.A(new_n875), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n384), .A2(new_n273), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n385), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n396), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n419), .B1(new_n889), .B2(new_n667), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n408), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n414), .A2(new_n416), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n667), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n398), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n889), .A2(new_n667), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n422), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n872), .A2(new_n885), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n660), .A2(new_n895), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT103), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n871), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n824), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n903), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n884), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  INV_X1    g0711(.A(new_n905), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n894), .B1(new_n893), .B2(new_n896), .ZN(new_n914));
  AND4_X1   g0714(.A1(new_n894), .A2(new_n410), .A3(new_n896), .A4(new_n419), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT105), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n410), .A2(new_n896), .A3(new_n419), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n897), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n422), .A2(new_n398), .A3(new_n895), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT106), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT39), .B1(new_n901), .B2(new_n902), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n925), .A4(new_n926), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(new_n371), .A4(new_n677), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n906), .A2(new_n913), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n711), .B(new_n438), .C1(new_n716), .C2(KEYINPUT29), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n662), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(G330), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n924), .A2(new_n926), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n733), .A2(new_n827), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n884), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT40), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n884), .A2(new_n939), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n438), .A2(new_n733), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n937), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n936), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n206), .B2(new_n739), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n936), .A2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n870), .B1(new_n950), .B2(new_n951), .ZN(G367));
  OAI221_X1 g0752(.A(new_n809), .B1(new_n210), .B2(new_n309), .C1(new_n798), .C2(new_n237), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n742), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT111), .Z(new_n955));
  OAI221_X1 g0755(.A(new_n515), .B1(new_n748), .B2(new_n300), .C1(new_n754), .C2(new_n849), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n779), .B2(G283), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n957), .B1(new_n522), .B2(new_n772), .C1(new_n958), .C2(new_n762), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n792), .A2(G116), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT46), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(new_n961), .B1(new_n757), .B2(G294), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .C1(new_n769), .C2(new_n845), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n779), .A2(G50), .B1(new_n784), .B2(G137), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n250), .B2(new_n772), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n251), .B1(new_n752), .B2(new_n753), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n789), .A2(new_n389), .B1(new_n748), .B2(new_n332), .ZN(new_n967));
  INV_X1    g0767(.A(new_n754), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n966), .B(new_n967), .C1(G150), .C2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n838), .B2(new_n769), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n959), .A2(new_n963), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT47), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n746), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n955), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n700), .A2(new_n677), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n638), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n703), .B2(new_n976), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(new_n811), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n596), .B(new_n603), .C1(new_n586), .C2(new_n677), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n644), .A2(new_n669), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n680), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n510), .A2(new_n681), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n981), .B2(new_n982), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT42), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n603), .B1(new_n981), .B2(new_n502), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n677), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT42), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n986), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT107), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n984), .B1(new_n985), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n985), .B2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n981), .A2(new_n982), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n682), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT45), .Z(new_n1003));
  NAND2_X1  g0803(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n682), .B2(new_n1001), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT110), .Z(new_n1007));
  XNOR2_X1  g0807(.A(new_n1005), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n680), .B(new_n1009), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n987), .B1(new_n679), .B2(new_n681), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n675), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n736), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n736), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n685), .B(KEYINPUT41), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n741), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n980), .B1(new_n1000), .B2(new_n1018), .ZN(G387));
  OR2_X1    g0819(.A1(new_n679), .A2(new_n811), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n801), .A2(new_n687), .B1(G107), .B2(new_n210), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n234), .A2(new_n458), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n687), .ZN(new_n1023));
  AOI211_X1 g0823(.A(G45), .B(new_n1023), .C1(G68), .C2(G77), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n277), .A2(G50), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n798), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1021), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n809), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n742), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n779), .A2(G68), .B1(new_n782), .B2(G97), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n784), .A2(G150), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n770), .A2(G159), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n251), .B1(new_n752), .B2(new_n250), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n789), .A2(new_n277), .B1(new_n309), .B2(new_n748), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G50), .C2(new_n968), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n251), .B1(new_n784), .B2(G326), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n752), .A2(new_n443), .B1(new_n748), .B2(new_n851), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n968), .A2(G317), .B1(G311), .B2(new_n757), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n787), .B2(new_n769), .C1(new_n778), .C2(new_n849), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1038), .B1(new_n524), .B2(new_n772), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1037), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1030), .B1(new_n1048), .B2(new_n745), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1012), .A2(new_n741), .B1(new_n1020), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1013), .A2(new_n685), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n736), .A2(new_n1012), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(G393));
  NAND2_X1  g0853(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1014), .A2(new_n1054), .A3(new_n685), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1001), .A2(new_n811), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n797), .A2(new_n241), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n809), .C1(new_n522), .C2(new_n210), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n796), .B1(new_n1058), .B2(KEYINPUT113), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n769), .A2(new_n958), .B1(new_n845), .B2(new_n754), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n773), .B1(new_n779), .B2(G294), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n787), .B2(new_n762), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n748), .A2(new_n524), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n515), .B1(new_n752), .B2(new_n851), .C1(new_n849), .C2(new_n789), .ZN(new_n1066));
  OR4_X1    g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n560), .A2(new_n772), .B1(new_n762), .B2(new_n838), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n515), .B1(new_n792), .B2(G68), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n250), .B2(new_n748), .C1(new_n789), .C2(new_n202), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(new_n307), .C2(new_n779), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n769), .A2(new_n279), .B1(new_n389), .B2(new_n754), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1059), .B1(KEYINPUT113), .B2(new_n1058), .C1(new_n1075), .C2(new_n746), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1010), .B(KEYINPUT112), .Z(new_n1077));
  OAI221_X1 g0877(.A(new_n1055), .B1(new_n1056), .B2(new_n1076), .C1(new_n1077), .C2(new_n740), .ZN(G390));
  AOI22_X1  g0878(.A1(new_n779), .A2(G97), .B1(G107), .B2(new_n757), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n851), .B2(new_n769), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT118), .Z(new_n1081));
  NOR2_X1   g0881(.A1(new_n748), .A2(new_n250), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n515), .B1(new_n752), .B2(new_n560), .C1(new_n524), .C2(new_n754), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n332), .A2(new_n772), .B1(new_n762), .B2(new_n443), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n792), .A2(G150), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1086), .A2(KEYINPUT53), .B1(new_n837), .B2(new_n754), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n779), .B2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n789), .A2(new_n840), .B1(new_n748), .B2(new_n389), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(KEYINPUT53), .B2(new_n1086), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G125), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n251), .B1(new_n762), .B2(new_n1093), .C1(new_n202), .C2(new_n772), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT117), .Z(new_n1095));
  AOI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(G128), .C2(new_n770), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n745), .B1(new_n1085), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n796), .B1(new_n277), .B2(new_n831), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n930), .A2(new_n931), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n806), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n733), .A2(new_n827), .A3(G330), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n884), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n908), .A2(new_n884), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n371), .A2(new_n677), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1106), .A2(new_n1107), .B1(new_n930), .B2(new_n931), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n938), .A2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n907), .B1(new_n707), .B2(new_n819), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT115), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n907), .C1(new_n707), .C2(new_n819), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n884), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1105), .B1(new_n1108), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n872), .B2(new_n885), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1100), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n1115), .A3(new_n1104), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1101), .B1(new_n1121), .B2(new_n741), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1102), .B(new_n877), .C1(new_n883), .C2(new_n882), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1104), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n872), .B1(new_n1104), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n438), .A2(new_n734), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n934), .A2(new_n662), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT116), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT116), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n1121), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1117), .A2(new_n1130), .A3(new_n1120), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n685), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1122), .B1(new_n1135), .B2(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(new_n932), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n291), .A2(new_n296), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n285), .A2(new_n895), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1142), .B(new_n1143), .Z(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1144), .B(new_n1145), .Z(new_n1146));
  NAND3_X1  g0946(.A1(new_n945), .A2(G330), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1144), .B(new_n1145), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(KEYINPUT40), .A2(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n937), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1141), .A2(new_n913), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1149), .A2(new_n937), .A3(new_n1148), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1146), .B1(new_n945), .B2(G330), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n933), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1129), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1136), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1151), .A2(new_n1154), .B1(new_n1136), .B2(new_n1156), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT57), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n685), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n742), .B1(G50), .B2(new_n832), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n782), .A2(G58), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n851), .B2(new_n762), .C1(new_n778), .C2(new_n309), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n769), .A2(new_n524), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n251), .A2(G41), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n752), .B2(new_n250), .C1(new_n300), .C2(new_n754), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n789), .A2(new_n522), .B1(new_n748), .B2(new_n332), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1171), .A2(KEYINPUT58), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT58), .B2(new_n1171), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n784), .A2(G124), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G33), .B(G41), .C1(new_n782), .C2(G159), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n968), .A2(G128), .B1(new_n792), .B2(new_n1088), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n279), .B2(new_n748), .C1(new_n769), .C2(new_n1093), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n779), .A2(G137), .B1(G132), .B2(new_n757), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT119), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT119), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1178), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT59), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1175), .B(new_n1176), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1174), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1164), .B1(new_n1187), .B2(new_n745), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1146), .B2(new_n807), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1155), .B2(new_n741), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1163), .A2(new_n1191), .ZN(G375));
  AOI21_X1  g0992(.A(new_n1016), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1132), .A2(new_n1133), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n742), .B1(G68), .B2(new_n832), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT122), .Z(new_n1199));
  OAI22_X1  g0999(.A1(new_n789), .A2(new_n524), .B1(new_n748), .B2(new_n309), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n515), .B1(new_n752), .B2(new_n522), .C1(new_n851), .C2(new_n754), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G294), .C2(new_n770), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G77), .A2(new_n782), .B1(new_n784), .B2(G303), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n300), .C2(new_n778), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1165), .A2(new_n251), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT123), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n779), .A2(G150), .B1(new_n784), .B2(G128), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n748), .A2(new_n202), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n754), .A2(new_n840), .B1(new_n752), .B2(new_n389), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n757), .C2(new_n1088), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1207), .B(new_n1210), .C1(new_n837), .C2(new_n769), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1199), .B1(new_n1212), .B2(new_n745), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n884), .B2(new_n807), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n740), .B(KEYINPUT121), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1127), .B2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT124), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1196), .A2(new_n1197), .A3(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT125), .Z(G381));
  OR2_X1    g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  OR4_X1    g1020(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1220), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G378), .A2(new_n1221), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1022(.A(G378), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n668), .A2(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(G375), .C2(new_n1226), .ZN(G409));
  XNOR2_X1  g1027(.A(G393), .B(new_n813), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(G390), .B(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(G387), .Z(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT61), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT127), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT60), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1130), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n685), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1217), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n830), .A3(new_n858), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(G384), .A3(new_n1217), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1225), .A2(G2897), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1161), .A2(new_n1017), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1215), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1190), .B1(new_n1155), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G378), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n685), .B1(new_n1161), .B2(KEYINPUT57), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1155), .A2(KEYINPUT57), .A3(new_n1157), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1191), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1163), .A2(new_n1252), .A3(G378), .A4(new_n1191), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1247), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1243), .B1(new_n1254), .B2(new_n1225), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1254), .A2(new_n1225), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1232), .B(new_n1255), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1247), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1256), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1224), .A3(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1231), .B1(new_n1259), .B2(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1255), .A2(new_n1232), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1257), .A2(KEYINPUT63), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1230), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1271), .ZN(G405));
  INV_X1    g1072(.A(G375), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1260), .B1(G378), .B2(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1274), .A2(new_n1263), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1263), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1230), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1231), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G402));
endmodule


