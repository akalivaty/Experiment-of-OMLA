//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n456));
  XOR2_X1   g031(.A(new_n455), .B(new_n456), .Z(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g035(.A(G261), .ZN(G325));
  INV_X1    g036(.A(new_n457), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2106), .ZN(new_n463));
  INV_X1    g038(.A(new_n458), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G567), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(G137), .A3(new_n468), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n479));
  INV_X1    g054(.A(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT3), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(new_n468), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n479), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n481), .A2(new_n483), .A3(G126), .A4(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n481), .A2(new_n483), .A3(G138), .A4(new_n468), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n469), .A2(new_n499), .A3(G138), .A4(new_n468), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(G543), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT72), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT70), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n510), .A2(new_n511), .A3(new_n517), .A4(new_n502), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n505), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n510), .A2(G62), .A3(new_n511), .A4(new_n517), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n518), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n504), .A2(G51), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n510), .A2(new_n511), .A3(new_n517), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n527), .A2(new_n534), .ZN(G168));
  NAND4_X1  g110(.A1(new_n510), .A2(G64), .A3(new_n511), .A4(new_n517), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n521), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G52), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n504), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n540), .B(new_n544), .C1(new_n518), .C2(new_n541), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n538), .B1(new_n543), .B2(new_n545), .ZN(G171));
  AND3_X1   g121(.A1(new_n510), .A2(new_n511), .A3(new_n517), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n521), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n504), .A2(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n518), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n504), .A2(G53), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n526), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n510), .A2(G65), .A3(new_n511), .A4(new_n517), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n568), .B2(G651), .ZN(new_n569));
  AOI211_X1 g144(.A(KEYINPUT76), .B(new_n521), .C1(new_n566), .C2(new_n567), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n563), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  NOR2_X1   g151(.A1(G171), .A2(KEYINPUT78), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  AOI211_X1 g153(.A(new_n578), .B(new_n538), .C1(new_n543), .C2(new_n545), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G301));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n547), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n526), .A2(G87), .B1(G49), .B2(new_n504), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n532), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n504), .A2(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(G651), .B2(new_n592), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n547), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n521), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT81), .B(G47), .Z(new_n605));
  OAI22_X1  g180(.A1(new_n518), .A2(new_n604), .B1(new_n503), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n532), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n504), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT10), .B1(new_n518), .B2(new_n613), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n518), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n580), .B2(new_n617), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(new_n580), .B2(new_n617), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n575), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n575), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT82), .B(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(G860), .B2(new_n625), .ZN(G148));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n485), .A2(G135), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT83), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n487), .A2(G123), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2100), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT84), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n658), .B2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n645), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n644), .A3(new_n663), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n668), .A3(G14), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT86), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n671));
  NAND4_X1  g246(.A1(new_n666), .A2(new_n668), .A3(new_n671), .A4(G14), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n675), .B1(new_n679), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT17), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n677), .A2(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n679), .B(new_n684), .C1(new_n682), .C2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n681), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n702), .B(new_n703), .C1(new_n701), .C2(new_n700), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(G229));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G35), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n489), .B2(G29), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n717), .A2(new_n718), .A3(G2090), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT97), .ZN(new_n720));
  OAI21_X1  g295(.A(G2090), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  NAND2_X1  g296(.A1(G164), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G27), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT30), .B(G28), .Z(new_n727));
  OAI211_X1 g302(.A(new_n725), .B(new_n726), .C1(G29), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n485), .A2(G139), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n468), .C2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G33), .B(new_n733), .S(G29), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2072), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n485), .A2(G141), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n487), .A2(G129), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT26), .Z(new_n740));
  NAND4_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G32), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(KEYINPUT27), .B(G1996), .Z(new_n743));
  OAI21_X1  g318(.A(new_n735), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT24), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n745), .B2(KEYINPUT24), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  AOI22_X1  g323(.A1(G160), .A2(G29), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n734), .A2(G2072), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n728), .A2(new_n744), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G16), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n755), .ZN(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n554), .B2(G16), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n759), .A2(new_n760), .B1(G1341), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n720), .A2(new_n721), .A3(new_n754), .A4(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n632), .A2(new_n713), .A3(new_n636), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT31), .B(G11), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n713), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT93), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n487), .A2(G128), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n485), .A2(G140), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n468), .A2(G116), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n769), .B1(new_n778), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2067), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n755), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n755), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT95), .Z(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n742), .A2(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n785), .A2(new_n786), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n755), .A2(KEYINPUT23), .A3(G20), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n793));
  INV_X1    g368(.A(G20), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G16), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n795), .C1(new_n575), .C2(new_n755), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n782), .A2(new_n790), .A3(new_n791), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n755), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n624), .B2(new_n755), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1348), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n762), .A2(G1341), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n755), .B1(new_n597), .B2(new_n600), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n755), .A2(G6), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n805), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(G16), .A2(G23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G288), .B2(new_n755), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G166), .A2(new_n755), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n755), .A2(G22), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n817), .A2(G1971), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(G1971), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n812), .B(new_n814), .C1(G288), .C2(new_n755), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n816), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n822), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n826), .A2(new_n824), .A3(new_n809), .A4(new_n810), .ZN(new_n827));
  AOI22_X1  g402(.A1(G119), .A2(new_n487), .B1(new_n485), .B2(G131), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n829));
  NOR2_X1   g404(.A1(G95), .A2(G2105), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT90), .Z(new_n831));
  OAI21_X1  g406(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G25), .B(new_n832), .S(G29), .Z(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT35), .B(G1991), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  NOR2_X1   g410(.A1(G16), .A2(G24), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n607), .B2(G16), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(G1986), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(G1986), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n827), .A2(new_n835), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT91), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n823), .A2(new_n824), .B1(G1986), .B2(new_n837), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT91), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n835), .A4(new_n838), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n825), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g422(.A(KEYINPUT36), .B(new_n825), .C1(new_n841), .C2(new_n844), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n804), .B1(new_n847), .B2(new_n848), .ZN(G150));
  NAND2_X1  g424(.A1(G150), .A2(KEYINPUT98), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n804), .B(new_n851), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G311));
  AOI22_X1  g428(.A1(new_n526), .A2(G93), .B1(G55), .B2(new_n504), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n532), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G651), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n554), .A2(new_n859), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n858), .B(new_n854), .C1(new_n550), .C2(new_n553), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT39), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n624), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n869), .B2(G860), .ZN(G145));
  XNOR2_X1  g445(.A(new_n778), .B(new_n733), .ZN(new_n871));
  INV_X1    g446(.A(G164), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n832), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n489), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n637), .ZN(new_n877));
  INV_X1    g452(.A(new_n640), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(G130), .A2(new_n487), .B1(new_n485), .B2(G142), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT100), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(KEYINPUT100), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n887), .B(new_n888), .C1(G118), .C2(new_n468), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(new_n741), .Z(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT101), .Z(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n882), .A2(new_n892), .A3(new_n883), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n573), .A2(new_n574), .A3(new_n616), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n569), .A2(new_n570), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(KEYINPUT77), .A3(new_n563), .A4(new_n564), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n571), .A2(new_n572), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n624), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n865), .B(new_n627), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT41), .B1(new_n900), .B2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n616), .B1(new_n573), .B2(new_n574), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n902), .A2(new_n903), .A3(new_n624), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G288), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G290), .ZN(new_n915));
  NAND2_X1  g490(.A1(G288), .A2(new_n607), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G305), .A2(G166), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n597), .A2(new_n600), .A3(G303), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n915), .A2(new_n918), .A3(new_n919), .A4(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(KEYINPUT42), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n907), .B(new_n913), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n907), .A2(new_n913), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(KEYINPUT102), .A3(new_n926), .A4(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(KEYINPUT103), .A3(G868), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n859), .B2(new_n617), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n933), .B2(G868), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n899), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n933), .A2(G868), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT104), .B(new_n934), .C1(new_n940), .C2(new_n937), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(G295));
  OAI21_X1  g517(.A(new_n934), .B1(new_n940), .B2(new_n937), .ZN(G331));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n908), .A2(new_n912), .ZN(new_n945));
  OAI21_X1  g520(.A(G168), .B1(new_n577), .B2(new_n579), .ZN(new_n946));
  NAND2_X1  g521(.A1(G286), .A2(G171), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n865), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n863), .A2(new_n864), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n946), .A2(new_n950), .A3(KEYINPUT105), .A4(new_n947), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n909), .A2(new_n911), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n950), .B1(new_n946), .B2(new_n947), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n923), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n944), .B1(new_n962), .B2(G37), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n953), .A2(new_n961), .A3(new_n923), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n945), .A2(new_n952), .B1(new_n957), .B2(new_n960), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT106), .B(new_n895), .C1(new_n965), .C2(new_n923), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n967), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n905), .A2(new_n949), .A3(new_n951), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n957), .A2(new_n949), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n912), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n909), .A2(KEYINPUT107), .A3(new_n910), .A4(new_n911), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n908), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n895), .B(new_n964), .C1(new_n976), .C2(new_n923), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n969), .B1(new_n977), .B2(KEYINPUT43), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT108), .B1(new_n967), .B2(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n968), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n969), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n980), .A2(new_n985), .ZN(G397));
  NAND2_X1  g561(.A1(new_n498), .A2(new_n500), .ZN(new_n987));
  INV_X1    g562(.A(new_n496), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT109), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G125), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n471), .B1(new_n484), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G2105), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(G40), .A3(new_n474), .A4(new_n473), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n999));
  OR3_X1    g574(.A1(new_n998), .A2(new_n999), .A3(G1996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n778), .A2(G2067), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n780), .A3(new_n777), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n1003), .B2(new_n741), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n999), .B1(new_n998), .B2(G1996), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1000), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  AND2_X1   g582(.A1(new_n997), .A2(new_n1003), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n741), .B(G1996), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1010), .B(new_n1011), .C1(new_n997), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n832), .A2(new_n834), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n998), .B1(new_n1015), .B2(new_n1002), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n832), .A2(new_n834), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n997), .B1(new_n1017), .B2(new_n1014), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(G290), .A2(G1986), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n998), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1007), .B(new_n1016), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n593), .B2(new_n596), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n598), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1025), .B(new_n1027), .C1(new_n1029), .C2(KEYINPUT49), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n472), .A2(new_n475), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n989), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G288), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n586), .A2(G1976), .A3(new_n587), .A4(new_n588), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1036), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1036), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n520), .B2(new_n524), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT55), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1048));
  INV_X1    g623(.A(new_n991), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(new_n1034), .C1(new_n989), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n996), .B1(new_n989), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n989), .B2(new_n1053), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1052), .B1(G2090), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1047), .A2(new_n1059), .A3(G8), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1054), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1052), .B1(G2090), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1047), .B1(new_n1064), .B2(G8), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1045), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1054), .A2(new_n1055), .A3(new_n751), .A4(new_n1057), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1034), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n989), .B2(new_n1049), .ZN(new_n1070));
  NOR4_X1   g645(.A1(G164), .A2(KEYINPUT114), .A3(G1384), .A4(new_n991), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(G168), .B(new_n1067), .C1(new_n1072), .C2(G1966), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(KEYINPUT122), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1067), .B1(new_n1072), .B2(G1966), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(G8), .A3(G286), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1074), .A2(new_n1081), .A3(new_n1075), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1058), .A2(KEYINPUT119), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1054), .A2(new_n1055), .A3(new_n1085), .A4(new_n1057), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n786), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1050), .B2(G2078), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1072), .A2(KEYINPUT53), .A3(new_n724), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n580), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1088), .A2(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n992), .A2(new_n1034), .A3(new_n1048), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1087), .A2(new_n1094), .A3(new_n1089), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n580), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(G171), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(KEYINPUT54), .C1(new_n580), .C2(new_n1091), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n1066), .A2(new_n1083), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1050), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1102), .A2(new_n1103), .B1(new_n1063), .B2(new_n797), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n563), .A3(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n571), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT118), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1116), .B(new_n1113), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1104), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1115), .A2(new_n1117), .A3(new_n1104), .ZN(new_n1119));
  INV_X1    g694(.A(G1348), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1084), .A2(new_n1120), .A3(new_n1086), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1034), .A2(new_n989), .A3(new_n780), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n616), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1118), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT121), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n1118), .C1(new_n1119), .C2(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1116), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1111), .A2(KEYINPUT118), .A3(new_n1114), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1104), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1135), .A2(new_n1118), .A3(KEYINPUT61), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT61), .B1(new_n1135), .B2(new_n1118), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n624), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n1139), .B2(new_n1123), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1035), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1050), .B2(G1996), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n554), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT59), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1140), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1136), .A2(new_n1137), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1101), .B1(new_n1130), .B2(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1045), .A2(new_n1060), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1037), .A2(new_n1038), .A3(new_n914), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n593), .A2(G1981), .A3(new_n596), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1036), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1079), .A2(G8), .A3(G168), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1079), .A2(KEYINPUT115), .A3(G8), .A4(G168), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n1066), .B2(new_n1158), .ZN(new_n1159));
  AND4_X1   g734(.A1(new_n1060), .A2(new_n1037), .A3(new_n1044), .A4(new_n1042), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1059), .A2(G8), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1047), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1160), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1150), .B(new_n1153), .C1(new_n1159), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1083), .A2(new_n1167), .A3(KEYINPUT62), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1083), .B2(KEYINPUT62), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1066), .A2(new_n580), .A3(new_n1091), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1166), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1149), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1020), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n997), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1019), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1182), .B(new_n1179), .C1(new_n1149), .C2(new_n1174), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1024), .B1(new_n1181), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n982), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n897), .A2(new_n711), .ZN(new_n1188));
  INV_X1    g762(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n466), .B1(new_n670), .B2(new_n672), .ZN(new_n1190));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1191));
  AND3_X1   g765(.A1(new_n1190), .A2(new_n1191), .A3(new_n690), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1190), .B2(new_n690), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1186), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1190), .A2(new_n690), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1196), .A2(KEYINPUT126), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1190), .A2(new_n1191), .A3(new_n690), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1188), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n984), .A2(new_n1199), .A3(KEYINPUT127), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1195), .A2(new_n1200), .ZN(G308));
  NAND2_X1  g775(.A1(new_n984), .A2(new_n1199), .ZN(G225));
endmodule


