//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n207), .B2(KEYINPUT87), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209));
  NOR2_X1   g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(new_n204), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n208), .A2(new_n211), .B1(new_n205), .B2(new_n206), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  OR3_X1    g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT15), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n207), .A2(new_n203), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT15), .B1(new_n213), .B2(new_n215), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n220), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(G1gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT16), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G1gat), .B2(new_n227), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(G8gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT90), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n220), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT90), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n226), .A2(new_n238), .A3(new_n233), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n202), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n226), .B2(new_n233), .ZN(new_n243));
  AOI211_X1 g042(.A(KEYINPUT90), .B(new_n232), .C1(new_n221), .C2(new_n225), .ZN(new_n244));
  INV_X1    g043(.A(new_n237), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n246), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(new_n236), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n241), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n220), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT13), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n242), .A2(new_n247), .A3(new_n248), .A4(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n256));
  XOR2_X1   g055(.A(G113gat), .B(G141gat), .Z(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G169gat), .B(G197gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT12), .Z(new_n262));
  AND3_X1   g061(.A1(new_n255), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n256), .B1(new_n255), .B2(new_n262), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n242), .A2(new_n247), .A3(new_n254), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n240), .A2(KEYINPUT93), .A3(new_n241), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT93), .B1(new_n240), .B2(new_n241), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  OAI22_X1  g068(.A1(new_n263), .A2(new_n264), .B1(new_n269), .B2(new_n262), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT23), .B(new_n273), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT66), .B(G176gat), .Z(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT23), .A4(new_n273), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT23), .B1(new_n273), .B2(new_n276), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G169gat), .B2(G176gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n287), .B2(KEYINPUT24), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT65), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n279), .A2(new_n282), .A3(new_n284), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n288), .A2(new_n290), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n273), .A2(new_n276), .A3(KEYINPUT23), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n284), .A4(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n298), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT69), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT69), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n305), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315));
  AOI21_X1  g114(.A(G190gat), .B1(new_n307), .B2(KEYINPUT69), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n316), .B(KEYINPUT70), .C1(KEYINPUT69), .C2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(KEYINPUT28), .A3(new_n309), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT26), .B1(new_n273), .B2(new_n276), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n273), .B2(new_n276), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n273), .A2(new_n276), .A3(KEYINPUT26), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n321), .A2(new_n323), .A3(new_n324), .A4(new_n286), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n272), .B1(new_n304), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G226gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n295), .A2(new_n297), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT68), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n302), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n325), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT22), .ZN(new_n338));
  NAND2_X1  g137(.A1(G211gat), .A2(G218gat), .ZN(new_n339));
  INV_X1    g138(.A(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(G218gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n334), .A2(new_n325), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n330), .A2(KEYINPUT29), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n349), .A2(new_n328), .A3(new_n329), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n335), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n352), .B1(new_n355), .B2(new_n348), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT37), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n351), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n347), .ZN(new_n360));
  INV_X1    g159(.A(new_n335), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT74), .B1(new_n334), .B2(new_n325), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n353), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n360), .B(KEYINPUT37), .C1(new_n365), .C2(new_n347), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  INV_X1    g166(.A(G64gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G92gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n358), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT38), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT37), .B(new_n352), .C1(new_n355), .C2(new_n348), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n375), .A2(KEYINPUT38), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n358), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  AND2_X1   g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G141gat), .B(G148gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(G155gat), .B2(G162gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G141gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G148gat), .ZN(new_n388));
  INV_X1    g187(.A(G148gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G141gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G155gat), .B(G162gat), .ZN(new_n392));
  INV_X1    g191(.A(G155gat), .ZN(new_n393));
  INV_X1    g192(.A(G162gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT2), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT3), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n386), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G113gat), .B(G120gat), .ZN(new_n401));
  OAI21_X1  g200(.A(G127gat), .B1(new_n401), .B2(KEYINPUT1), .ZN(new_n402));
  INV_X1    g201(.A(G120gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(G113gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G120gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n408));
  INV_X1    g207(.A(G127gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(new_n410), .A3(G134gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(G134gat), .B1(new_n402), .B2(new_n410), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n398), .B(new_n400), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G134gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n407), .B2(new_n408), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT1), .B(G127gat), .C1(new_n404), .C2(new_n406), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n386), .A2(new_n396), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n411), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT75), .B1(new_n420), .B2(KEYINPUT4), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT76), .A4(new_n411), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT4), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n379), .B(new_n414), .C1(new_n424), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n411), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n397), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  INV_X1    g232(.A(new_n379), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n426), .B2(new_n427), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n412), .A2(new_n413), .A3(new_n397), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n414), .B2(KEYINPUT4), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n379), .A2(new_n430), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G1gat), .B(G29gat), .Z(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454));
  INV_X1    g253(.A(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n434), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n420), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(new_n421), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n426), .A2(new_n427), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n437), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n434), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n462), .B2(new_n414), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT83), .B1(new_n463), .B2(new_n442), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n436), .A2(new_n465), .A3(new_n443), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n455), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n451), .B1(new_n444), .B2(new_n449), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n454), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n465), .B1(new_n436), .B2(new_n443), .ZN(new_n470));
  AOI211_X1 g269(.A(KEYINPUT83), .B(new_n442), .C1(new_n429), .C2(new_n435), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n449), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n463), .A2(new_n442), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT6), .B1(new_n473), .B2(new_n455), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT85), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n371), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n356), .B2(KEYINPUT38), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n378), .A2(new_n453), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n399), .B1(new_n347), .B2(KEYINPUT29), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n397), .ZN(new_n481));
  INV_X1    g280(.A(G228gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n329), .ZN(new_n483));
  INV_X1    g282(.A(new_n400), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n347), .B1(new_n484), .B2(KEYINPUT29), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n343), .A2(KEYINPUT78), .A3(new_n346), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n397), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n398), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT79), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(KEYINPUT79), .A3(new_n398), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n485), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n483), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT80), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n487), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G22gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G78gat), .B(G106gat), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT31), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n502), .A2(KEYINPUT81), .A3(new_n503), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT81), .B1(new_n502), .B2(new_n503), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n502), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT82), .B1(new_n514), .B2(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT82), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n502), .A2(new_n516), .A3(new_n503), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n510), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n356), .A2(KEYINPUT30), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(new_n352), .C1(new_n355), .C2(new_n348), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(new_n477), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n356), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n438), .A2(new_n440), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n525), .A2(KEYINPUT39), .A3(new_n379), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n449), .B1(KEYINPUT84), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(new_n379), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT39), .B1(new_n433), .B2(new_n434), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n526), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n527), .A2(KEYINPUT84), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n523), .A2(new_n524), .A3(new_n533), .A4(new_n472), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n479), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT64), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n431), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n334), .A2(new_n541), .A3(new_n325), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n334), .B2(new_n325), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT32), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G43gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(G71gat), .B(G99gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n544), .B(KEYINPUT32), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT71), .B1(new_n542), .B2(new_n543), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n349), .A2(new_n431), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n334), .A2(new_n541), .A3(new_n325), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n559), .A3(new_n538), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT34), .ZN(new_n561));
  OR4_X1    g360(.A1(KEYINPUT34), .A2(new_n542), .A3(new_n543), .A4(new_n540), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n551), .A2(new_n561), .A3(new_n553), .A4(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT73), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n569), .B(KEYINPUT36), .C1(new_n564), .C2(new_n565), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n563), .A3(KEYINPUT72), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n567), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n519), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n474), .A2(new_n450), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n453), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n523), .ZN(new_n581));
  INV_X1    g380(.A(new_n524), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n537), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n573), .A2(new_n574), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n519), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT35), .B1(new_n587), .B2(new_n583), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n581), .A2(new_n582), .ZN(new_n589));
  INV_X1    g388(.A(new_n566), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n469), .A2(new_n453), .A3(new_n475), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n519), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n588), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n271), .B1(new_n585), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT94), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n368), .A2(G57gat), .ZN(new_n602));
  INV_X1    g401(.A(G57gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(G64gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n604), .B(KEYINPUT95), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n601), .B(new_n596), .C1(new_n607), .C2(new_n602), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n232), .B1(new_n609), .B2(KEYINPUT21), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G183gat), .ZN(new_n611));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT96), .B(G211gat), .Z(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n613), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(G92gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(G85gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(KEYINPUT8), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT7), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT97), .B1(G85gat), .B2(G92gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n627), .ZN(new_n634));
  NOR2_X1   g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n633), .A2(KEYINPUT99), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n628), .B(new_n632), .C1(new_n634), .C2(new_n635), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(KEYINPUT99), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n226), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n637), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n642), .A2(new_n220), .B1(KEYINPUT100), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n646));
  NAND2_X1  g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n641), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G134gat), .B(G162gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n646), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n609), .A2(new_n638), .A3(new_n639), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n642), .B2(new_n609), .ZN(new_n659));
  INV_X1    g458(.A(G230gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n329), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT101), .Z(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n664), .B(new_n658), .C1(new_n642), .C2(new_n609), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n642), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n276), .ZN(new_n671));
  INV_X1    g470(.A(G204gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n663), .A2(new_n675), .A3(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n624), .A2(new_n657), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n595), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n580), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n589), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT103), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT105), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n686), .B1(new_n688), .B2(KEYINPUT104), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(KEYINPUT104), .B2(new_n688), .ZN(new_n692));
  OAI22_X1  g491(.A1(new_n685), .A2(new_n692), .B1(new_n686), .B2(G8gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(G1325gat));
  AOI21_X1  g493(.A(G15gat), .B1(new_n681), .B2(new_n590), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n575), .A2(new_n568), .A3(new_n570), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n681), .B2(new_n697), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n578), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  XNOR2_X1  g500(.A(new_n677), .B(KEYINPUT106), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n271), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  INV_X1    g505(.A(new_n657), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n706), .B(new_n707), .C1(new_n585), .C2(new_n594), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n372), .A2(new_n373), .B1(new_n376), .B2(new_n358), .ZN(new_n710));
  INV_X1    g509(.A(new_n478), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n591), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n584), .B1(new_n712), .B2(new_n535), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n713), .B2(new_n696), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n537), .A2(new_n577), .A3(KEYINPUT107), .A4(new_n584), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n594), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n657), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n705), .B(new_n708), .C1(new_n706), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n624), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n580), .ZN(new_n720));
  INV_X1    g519(.A(new_n624), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n677), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n595), .A2(new_n657), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n205), .A3(new_n682), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n720), .A2(new_n726), .ZN(G1328gat));
  INV_X1    g526(.A(new_n589), .ZN(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n719), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n723), .A2(G36gat), .A3(new_n728), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT46), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1329gat));
  AOI21_X1  g531(.A(new_n708), .B1(new_n717), .B2(new_n706), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(new_n696), .A3(new_n624), .A4(new_n704), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n736));
  INV_X1    g535(.A(G43gat), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n724), .A2(KEYINPUT108), .A3(new_n737), .A4(new_n590), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n595), .A2(new_n590), .A3(new_n657), .A4(new_n722), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(G43gat), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n736), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n735), .B(new_n742), .C1(KEYINPUT109), .C2(KEYINPUT47), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1330gat));
  NAND4_X1  g546(.A1(new_n718), .A2(G50gat), .A3(new_n578), .A4(new_n624), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n507), .B1(new_n723), .B2(new_n519), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1331gat));
  AND3_X1   g552(.A1(new_n716), .A2(new_n721), .A3(new_n707), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n703), .A2(new_n271), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n580), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n603), .ZN(G1332gat));
  XOR2_X1   g558(.A(new_n589), .B(KEYINPUT111), .Z(new_n760));
  NAND3_X1  g559(.A1(new_n754), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT49), .B(G64gat), .Z(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n761), .B2(new_n763), .ZN(G1333gat));
  XOR2_X1   g563(.A(new_n566), .B(KEYINPUT112), .Z(new_n765));
  AND3_X1   g564(.A1(new_n754), .A2(new_n756), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n696), .A2(G71gat), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n766), .A2(G71gat), .B1(new_n757), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g568(.A1(new_n757), .A2(new_n519), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(new_n600), .ZN(G1335gat));
  NAND2_X1  g570(.A1(new_n271), .A2(new_n624), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n677), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n774), .B(new_n708), .C1(new_n717), .C2(new_n706), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n580), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n716), .A2(new_n657), .A3(new_n773), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n716), .A2(KEYINPUT51), .A3(new_n657), .A4(new_n773), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n677), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n783), .A2(G85gat), .A3(new_n580), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT113), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n777), .A2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(new_n760), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n625), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n780), .B2(new_n781), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n702), .A2(G92gat), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n589), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n794), .A2(new_n625), .B1(new_n790), .B2(new_n791), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n776), .B2(new_n577), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n783), .A2(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n590), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1338gat));
  INV_X1    g600(.A(G106gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n775), .B2(new_n578), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n702), .A2(G106gat), .A3(new_n519), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT53), .B1(new_n782), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n805), .B(KEYINPUT114), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT115), .B1(new_n782), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n811), .B(new_n808), .C1(new_n780), .C2(new_n781), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n803), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n807), .B1(new_n813), .B2(new_n814), .ZN(G1339gat));
  NAND4_X1  g614(.A1(new_n242), .A2(new_n247), .A3(new_n266), .A4(new_n254), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n267), .A3(new_n262), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n246), .A2(new_n236), .B1(new_n251), .B2(new_n253), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n261), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n665), .A2(new_n661), .A3(new_n666), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n668), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n673), .B1(new_n668), .B2(KEYINPUT54), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n825), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n828), .A3(new_n676), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n820), .A2(new_n657), .A3(new_n830), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n270), .A2(new_n830), .B1(new_n820), .B2(new_n677), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n657), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n624), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n678), .A2(new_n271), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n587), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n682), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n835), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n833), .B2(new_n624), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n580), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT117), .A3(new_n837), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n760), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n405), .A3(new_n270), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n842), .A2(new_n578), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n760), .A2(new_n580), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n590), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT116), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n847), .A2(new_n851), .A3(new_n590), .A4(new_n848), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n850), .A2(new_n270), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n846), .B1(new_n853), .B2(new_n405), .ZN(G1340gat));
  NAND3_X1  g653(.A1(new_n845), .A2(new_n403), .A3(new_n677), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n850), .A2(new_n703), .A3(new_n852), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n403), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n845), .A2(KEYINPUT118), .A3(new_n721), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT117), .B1(new_n843), .B2(new_n837), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n842), .A2(new_n839), .A3(new_n580), .A4(new_n587), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n721), .B(new_n788), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n858), .A2(new_n863), .A3(new_n409), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n850), .A2(G127gat), .A3(new_n721), .A4(new_n852), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(G1342gat));
  NOR2_X1   g665(.A1(new_n589), .A2(new_n707), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n415), .B(new_n867), .C1(new_n859), .C2(new_n860), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(KEYINPUT120), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(KEYINPUT120), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n657), .A3(new_n852), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT119), .A3(G134gat), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n874), .B2(G134gat), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n871), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(G1343gat));
  NOR4_X1   g676(.A1(new_n842), .A2(new_n580), .A3(new_n696), .A4(new_n519), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n788), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n387), .B1(new_n879), .B2(new_n271), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n519), .B1(new_n834), .B2(new_n835), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT121), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n829), .B(KEYINPUT122), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n270), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n820), .A2(new_n677), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n657), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n831), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n624), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n835), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(KEYINPUT57), .A3(new_n578), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n891), .B(new_n892), .C1(new_n842), .C2(new_n519), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n882), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n760), .A2(new_n580), .A3(new_n696), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n270), .A2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n880), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT58), .B(new_n880), .C1(new_n896), .C2(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1344gat));
  NAND4_X1  g701(.A1(new_n878), .A2(new_n389), .A3(new_n677), .A4(new_n788), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n894), .A2(new_n677), .A3(new_n895), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(G148gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n679), .A2(new_n271), .A3(new_n680), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n888), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n578), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n836), .A2(new_n578), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n909), .A2(new_n911), .A3(new_n677), .A4(new_n895), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n905), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n903), .B1(new_n906), .B2(new_n913), .ZN(G1345gat));
  NAND2_X1  g713(.A1(new_n721), .A2(G155gat), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT123), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n895), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n393), .B1(new_n879), .B2(new_n624), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n896), .B2(new_n707), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n878), .A2(new_n394), .A3(new_n867), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n728), .A2(new_n682), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n836), .A2(new_n519), .A3(new_n765), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n271), .ZN(new_n925));
  NOR4_X1   g724(.A1(new_n842), .A2(new_n682), .A3(new_n587), .A4(new_n788), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n273), .A3(new_n270), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1348gat));
  NOR3_X1   g727(.A1(new_n924), .A2(new_n280), .A3(new_n702), .ZN(new_n929));
  AOI21_X1  g728(.A(G176gat), .B1(new_n926), .B2(new_n677), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n924), .A2(new_n932), .A3(new_n624), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n924), .B2(new_n624), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(G183gat), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n926), .A2(new_n317), .A3(new_n721), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  NAND4_X1  g740(.A1(new_n847), .A2(new_n657), .A3(new_n765), .A4(new_n923), .ZN(new_n942));
  NAND2_X1  g741(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(G190gat), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n309), .A3(new_n657), .ZN(new_n947));
  INV_X1    g746(.A(new_n945), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n942), .A2(G190gat), .A3(new_n948), .A4(new_n943), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n946), .A2(new_n949), .A3(new_n952), .A4(new_n947), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1351gat));
  NAND4_X1  g753(.A1(new_n909), .A2(new_n911), .A3(new_n577), .A4(new_n923), .ZN(new_n955));
  OAI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n271), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n842), .A2(new_n682), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n696), .A2(new_n519), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n760), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n271), .A2(G197gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n959), .A2(G204gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n677), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NOR4_X1   g764(.A1(new_n959), .A2(KEYINPUT127), .A3(G204gat), .A4(new_n783), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(KEYINPUT62), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n955), .B2(new_n702), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n964), .B2(new_n966), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(G1353gat));
  INV_X1    g771(.A(new_n959), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n340), .A3(new_n721), .ZN(new_n974));
  OAI211_X1 g773(.A(KEYINPUT63), .B(G211gat), .C1(new_n955), .C2(new_n624), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n908), .A2(new_n578), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n977), .A2(new_n577), .A3(new_n721), .A4(new_n923), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n974), .B1(new_n976), .B2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n955), .B2(new_n707), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n973), .A2(new_n341), .A3(new_n657), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


