//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT2), .B(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n201), .A3(KEYINPUT67), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n200), .A3(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n208), .A2(KEYINPUT64), .A3(G146), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT64), .B1(new_n208), .B2(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G146), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n211), .A2(new_n214), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT11), .B1(new_n218), .B2(G137), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G134), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT65), .B(G131), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n221), .B2(G134), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n218), .A3(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n223), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G131), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n226), .A2(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(new_n222), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n217), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n207), .A3(new_n215), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n208), .A2(G146), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n206), .B2(G143), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n208), .A2(KEYINPUT64), .A3(G146), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n237), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n232), .A2(new_n224), .A3(new_n233), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n218), .A2(G137), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n221), .A2(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n235), .A2(new_n236), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n236), .B1(new_n235), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n205), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT31), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n202), .A2(new_n204), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n235), .A2(new_n256), .A3(new_n251), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n254), .A2(new_n255), .A3(new_n257), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n207), .A2(new_n215), .A3(new_n212), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n212), .A2(new_n213), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n244), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(G131), .B1(new_n223), .B2(new_n229), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n247), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n205), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n266), .B1(new_n273), .B2(new_n257), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(new_n266), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT30), .B1(new_n267), .B2(new_n272), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n235), .A2(new_n236), .A3(new_n251), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n256), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n257), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n282), .A2(new_n283), .A3(new_n265), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n279), .B1(new_n284), .B2(new_n255), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n254), .A2(new_n257), .A3(new_n263), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n278), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G472), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT69), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(G472), .B2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n187), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT70), .B1(new_n288), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n273), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n283), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n275), .B(new_n263), .C1(new_n301), .C2(new_n266), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n254), .A2(new_n257), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n265), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n274), .A2(new_n276), .A3(new_n265), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n289), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n264), .A2(new_n277), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n286), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT68), .B1(new_n286), .B2(KEYINPUT31), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n297), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n296), .A2(new_n299), .A3(new_n310), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n294), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n309), .B1(new_n319), .B2(new_n187), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n299), .A4(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G217), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(G234), .B2(new_n290), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT73), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G137), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n195), .A2(G128), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n195), .A2(G128), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT24), .B(G110), .Z(new_n336));
  NAND3_X1  g150(.A1(new_n237), .A2(KEYINPUT23), .A3(G119), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(new_n334), .C1(new_n332), .C2(KEYINPUT23), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n335), .A2(new_n336), .B1(G110), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n340), .A2(KEYINPUT16), .A3(G140), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n206), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n335), .A2(new_n336), .ZN(new_n347));
  INV_X1    g161(.A(new_n341), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n340), .A2(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT16), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(new_n206), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n343), .A2(G146), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n338), .A2(KEYINPUT72), .A3(G110), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT72), .B1(new_n338), .B2(G110), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT74), .B(new_n346), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n206), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n344), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(new_n347), .C1(new_n359), .C2(new_n358), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT74), .B1(new_n365), .B2(new_n346), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n331), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n346), .B1(new_n357), .B2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT74), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n331), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n327), .B1(new_n372), .B2(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n369), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n361), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n370), .B1(new_n375), .B2(new_n331), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT25), .A3(new_n290), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n326), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n325), .A2(G902), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT75), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  OAI21_X1  g199(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT76), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT77), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  AOI21_X1  g212(.A(G101), .B1(new_n388), .B2(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n217), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(G104), .B1(new_n391), .B2(new_n393), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT78), .B1(new_n388), .B2(G107), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n390), .A3(G104), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G101), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(new_n400), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT10), .A3(new_n246), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n230), .A2(new_n234), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n239), .B1(new_n216), .B2(new_n245), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n400), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT10), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n405), .A2(new_n413), .A3(new_n414), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n416), .B1(new_n412), .B2(new_n246), .ZN(new_n420));
  INV_X1    g234(.A(new_n414), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(KEYINPUT12), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT12), .B1(new_n420), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G110), .B(G140), .ZN(new_n426));
  INV_X1    g240(.A(G227), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G953), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n426), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n405), .A2(new_n413), .A3(new_n418), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n421), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n425), .A2(new_n429), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G469), .B1(new_n435), .B2(G902), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  INV_X1    g251(.A(new_n424), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n431), .B1(new_n422), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n430), .B1(new_n434), .B2(new_n419), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n437), .B(new_n290), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n387), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n384), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n323), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n197), .A2(G119), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n188), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT5), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n450), .A2(new_n451), .B1(new_n193), .B2(new_n192), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n411), .A3(new_n400), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G104), .B2(new_n390), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT77), .B(G107), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n389), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n402), .B1(new_n458), .B2(new_n396), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n404), .A2(new_n202), .A3(new_n204), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n453), .B(new_n454), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n205), .A2(new_n401), .A3(new_n404), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n453), .A4(new_n454), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n453), .ZN(new_n470));
  INV_X1    g284(.A(new_n454), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n270), .A2(G125), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(G125), .B2(new_n246), .ZN(new_n477));
  INV_X1    g291(.A(G224), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n452), .A2(new_n411), .A3(new_n400), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n404), .A2(new_n202), .A3(new_n204), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n401), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n468), .A2(new_n472), .A3(KEYINPUT80), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n475), .A2(new_n480), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT6), .B1(new_n483), .B2(new_n454), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n467), .B2(new_n464), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n484), .B1(new_n491), .B2(KEYINPUT80), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT81), .A3(new_n480), .A4(new_n475), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n454), .B(KEYINPUT8), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n412), .A2(new_n452), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n481), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n477), .B1(new_n498), .B2(new_n479), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n477), .A2(new_n498), .A3(new_n479), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n502), .B2(new_n468), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G210), .B1(G237), .B2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n505), .A3(new_n503), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n447), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT83), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n258), .A2(new_n259), .A3(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n208), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n258), .A2(new_n259), .A3(G143), .A4(G214), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n225), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n513), .A3(new_n224), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n515), .A2(new_n516), .B1(G146), .B2(new_n343), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n342), .A2(KEYINPUT82), .A3(KEYINPUT19), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT19), .B1(new_n342), .B2(KEYINPUT82), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n206), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n231), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n514), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n352), .A2(G146), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n514), .A2(new_n523), .B1(new_n525), .B2(new_n345), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n517), .A2(new_n521), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n388), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n510), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n524), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n224), .B1(new_n512), .B2(new_n513), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n363), .A3(new_n344), .ZN(new_n534));
  INV_X1    g348(.A(new_n516), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n535), .A2(KEYINPUT17), .A3(new_n532), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n529), .B(new_n531), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n344), .B1(new_n535), .B2(new_n532), .ZN(new_n538));
  INV_X1    g352(.A(new_n520), .ZN(new_n539));
  AOI21_X1  g353(.A(G146), .B1(new_n539), .B2(new_n518), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n531), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n529), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(KEYINPUT83), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n530), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT84), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n530), .A2(new_n543), .A3(KEYINPUT84), .A4(new_n537), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT85), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n553));
  NOR3_X1   g367(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n531), .B1(new_n534), .B2(new_n536), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n542), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n537), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n290), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(G116), .B(G122), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n391), .A2(new_n393), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n564), .A2(KEYINPUT14), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n197), .A2(G122), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n390), .B1(new_n568), .B2(KEYINPUT14), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT86), .B1(new_n237), .B2(G143), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT86), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n208), .A3(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(G128), .B2(new_n208), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(G134), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(G134), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n570), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT87), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n570), .B(KEYINPUT87), .C1(new_n576), .C2(new_n577), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n577), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n564), .A2(new_n565), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT13), .B1(new_n571), .B2(new_n573), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT13), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n585), .B(new_n586), .C1(new_n237), .C2(G143), .ZN(new_n587));
  OAI221_X1 g401(.A(new_n583), .B1(new_n566), .B2(new_n584), .C1(new_n587), .C2(new_n218), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n385), .A2(new_n324), .A3(G953), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n582), .A2(new_n588), .A3(new_n590), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n290), .ZN(new_n595));
  INV_X1    g409(.A(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(KEYINPUT15), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n595), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(G902), .A3(G953), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT89), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT21), .B(G898), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT88), .B(G952), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(G953), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n602), .A2(new_n603), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT90), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n563), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n509), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n445), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n402), .ZN(G3));
  OAI21_X1  g426(.A(G472), .B1(new_n288), .B2(G902), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n383), .A2(new_n613), .A3(new_n442), .A4(new_n319), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT91), .Z(new_n615));
  NAND2_X1  g429(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT92), .B(KEYINPUT33), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n592), .A2(new_n593), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(G478), .A3(new_n290), .A4(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT93), .B(G478), .Z(new_n621));
  NAND2_X1  g435(.A1(new_n595), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n549), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT85), .B1(new_n549), .B2(KEYINPUT20), .ZN(new_n625));
  INV_X1    g439(.A(new_n555), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n623), .B1(new_n627), .B2(new_n561), .ZN(new_n628));
  INV_X1    g442(.A(new_n607), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n615), .A2(new_n509), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT94), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n546), .A2(new_n548), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n554), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n552), .A2(new_n553), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n595), .B(new_n597), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n562), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n509), .A2(KEYINPUT95), .A3(new_n607), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n505), .B1(new_n494), .B2(new_n503), .ZN(new_n644));
  INV_X1    g458(.A(new_n503), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n506), .B(new_n645), .C1(new_n489), .C2(new_n493), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n446), .B(new_n607), .C1(new_n644), .C2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n643), .B1(new_n647), .B2(new_n640), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n615), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n331), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n368), .B(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n380), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n378), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n443), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n613), .A2(new_n319), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n610), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT96), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n446), .B1(new_n644), .B2(new_n646), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n605), .A2(new_n600), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT97), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n602), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n638), .A2(new_n639), .A3(new_n562), .A4(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n664), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n657), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n318), .B2(new_n322), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n507), .A2(new_n508), .ZN(new_n675));
  INV_X1    g489(.A(new_n671), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT98), .A4(new_n446), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n672), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n672), .A2(new_n674), .A3(new_n677), .A4(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n675), .B(KEYINPUT38), .Z(new_n684));
  AND2_X1   g498(.A1(new_n299), .A2(new_n316), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n303), .A2(new_n263), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n301), .B2(new_n265), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n289), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n319), .B2(new_n187), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n599), .B1(new_n556), .B2(new_n562), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n446), .A3(new_n656), .A4(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n670), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n442), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT40), .Z(new_n698));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n556), .A2(new_n562), .B1(new_n622), .B2(new_n620), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n509), .A2(new_n701), .A3(new_n702), .A4(new_n670), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n623), .B(new_n670), .C1(new_n627), .C2(new_n561), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT101), .B1(new_n665), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n705), .A3(new_n674), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  OAI21_X1  g521(.A(new_n290), .B1(new_n439), .B2(new_n440), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n386), .A3(new_n441), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT102), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n712), .A3(new_n386), .A4(new_n441), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n711), .A2(new_n383), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n323), .A2(new_n630), .A3(new_n509), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND2_X1  g531(.A1(new_n323), .A2(new_n714), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n642), .B2(new_n648), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT103), .B(G116), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G18));
  INV_X1    g535(.A(new_n710), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n563), .A2(new_n608), .A3(new_n656), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n323), .A2(new_n509), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  AND3_X1   g539(.A1(new_n711), .A2(new_n607), .A3(new_n713), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n294), .B(KEYINPUT104), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n284), .A2(new_n255), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n278), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n613), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT105), .B1(new_n378), .B2(new_n382), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT25), .B1(new_n376), .B2(new_n290), .ZN(new_n732));
  AND4_X1   g546(.A1(KEYINPUT25), .A2(new_n367), .A3(new_n290), .A4(new_n371), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n325), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n381), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n509), .A2(new_n726), .A3(new_n691), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NAND2_X1  g554(.A1(new_n509), .A2(new_n722), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n656), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n730), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n704), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(new_n386), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n436), .B2(new_n441), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n644), .A2(new_n646), .A3(new_n447), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n323), .A3(new_n752), .A4(new_n383), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n296), .B(new_n310), .C1(new_n288), .C2(new_n298), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n702), .A2(new_n755), .A3(new_n670), .A4(new_n737), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n507), .A2(new_n446), .A3(new_n508), .A4(new_n749), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT42), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n753), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n754), .B1(new_n753), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND4_X1  g576(.A1(new_n751), .A2(new_n323), .A3(new_n383), .A4(new_n676), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NAND3_X1  g578(.A1(new_n556), .A2(new_n562), .A3(new_n623), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT43), .Z(new_n766));
  NOR2_X1   g580(.A1(new_n658), .A2(new_n656), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n644), .A2(new_n646), .A3(new_n447), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT110), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT110), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n775));
  OAI21_X1  g589(.A(G469), .B1(new_n435), .B2(KEYINPUT45), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT46), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n441), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n781), .B2(KEYINPUT107), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(KEYINPUT107), .B2(new_n781), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n386), .A3(new_n696), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(KEYINPUT108), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n773), .A2(new_n774), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  INV_X1    g604(.A(new_n770), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n791), .A2(new_n323), .A3(new_n383), .A4(new_n704), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT112), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n783), .A2(new_n386), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n783), .A2(new_n386), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(new_n796), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NAND2_X1  g615(.A1(new_n709), .A2(new_n441), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n447), .B(new_n387), .C1(new_n802), .C2(KEYINPUT49), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n804));
  INV_X1    g618(.A(new_n737), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n804), .A2(new_n690), .A3(new_n805), .A4(new_n765), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n684), .A2(new_n806), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n680), .A2(new_n681), .B1(new_n742), .B2(new_n745), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n656), .A2(new_n749), .A3(new_n670), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n690), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n691), .B(new_n446), .C1(new_n644), .C2(new_n646), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n810), .B1(new_n685), .B2(new_n689), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n509), .A2(new_n815), .A3(new_n816), .A4(new_n691), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n706), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n808), .A2(new_n809), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n809), .B1(new_n808), .B2(new_n819), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n562), .A2(new_n638), .A3(new_n599), .A4(new_n670), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n323), .A2(new_n657), .A3(new_n770), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n751), .A2(new_n745), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n763), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n763), .A2(new_n824), .A3(KEYINPUT113), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n556), .A2(new_n562), .A3(new_n639), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n614), .B1(new_n628), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n509), .A3(new_n607), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n715), .A2(new_n724), .A3(new_n739), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n610), .B1(new_n445), .B2(new_n659), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n834), .A2(new_n719), .A3(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n753), .A2(KEYINPUT53), .A3(new_n758), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n830), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n821), .A2(new_n822), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n840));
  NAND3_X1  g654(.A1(new_n830), .A2(new_n836), .A3(new_n761), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n682), .A2(new_n819), .A3(new_n746), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n830), .A2(new_n836), .A3(new_n761), .A4(KEYINPUT114), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n820), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(KEYINPUT54), .B(new_n839), .C1(new_n840), .C2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n840), .B2(new_n847), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n848), .B1(KEYINPUT54), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n684), .A2(new_n447), .A3(new_n722), .ZN(new_n853));
  INV_X1    g667(.A(new_n667), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n766), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n738), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT117), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n791), .A2(new_n710), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n744), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n690), .A2(new_n666), .A3(new_n384), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n563), .A2(new_n623), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n862), .A2(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n859), .A2(new_n860), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n859), .A2(KEYINPUT118), .A3(new_n860), .A4(new_n867), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n855), .A2(new_n738), .A3(new_n771), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n709), .A2(new_n387), .A3(new_n441), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n799), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n870), .A2(KEYINPUT51), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n859), .A2(new_n860), .A3(new_n867), .A4(new_n874), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n755), .A2(new_n737), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n862), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n865), .A2(new_n702), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n855), .A2(new_n742), .A3(new_n738), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n882), .A2(new_n605), .A3(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n875), .A2(new_n878), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(G952), .A2(G953), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT119), .B1(new_n852), .B2(new_n885), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n807), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n259), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n839), .B1(new_n847), .B2(new_n840), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n290), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(G210), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n492), .A2(new_n475), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n480), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n892), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n895), .B2(new_n899), .ZN(G51));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n439), .A2(new_n440), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n893), .B(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n778), .B(KEYINPUT57), .Z(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n893), .A2(new_n290), .A3(new_n777), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n902), .B(new_n892), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n847), .A2(new_n840), .ZN(new_n910));
  INV_X1    g724(.A(new_n839), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n906), .B1(new_n848), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n903), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT121), .B1(new_n915), .B2(new_n891), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n909), .A2(new_n916), .ZN(G54));
  AND3_X1   g731(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n892), .B1(new_n918), .B2(new_n636), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n636), .B2(new_n918), .ZN(G60));
  NAND2_X1  g734(.A1(new_n617), .A2(new_n619), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT122), .Z(new_n922));
  INV_X1    g736(.A(new_n852), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n905), .A2(new_n922), .A3(new_n925), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n892), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(new_n910), .A2(new_n911), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n654), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n930), .A2(new_n932), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n892), .B(new_n933), .C1(new_n934), .C2(new_n376), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n603), .B2(new_n478), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n836), .B2(G953), .ZN(new_n939));
  INV_X1    g753(.A(new_n896), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(G898), .B2(new_n259), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n939), .B(new_n942), .ZN(G69));
  NOR2_X1   g757(.A1(new_n519), .A2(new_n520), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n252), .A2(new_n253), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n697), .B(new_n791), .C1(new_n628), .C2(new_n831), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n383), .A3(new_n323), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n789), .A2(new_n800), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n808), .A2(new_n706), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n699), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n948), .B1(new_n956), .B2(G953), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n787), .A2(new_n509), .A3(new_n691), .A4(new_n879), .ZN(new_n958));
  AND4_X1   g772(.A1(new_n761), .A2(new_n958), .A3(new_n763), .A4(new_n800), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n789), .A2(KEYINPUT126), .A3(new_n952), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT126), .B1(new_n789), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n948), .A2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(G900), .B1(KEYINPUT127), .B2(G227), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n962), .A2(new_n963), .B1(G953), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n957), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n427), .B2(new_n668), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G72));
  OAI211_X1 g783(.A(new_n836), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  AOI211_X1 g786(.A(new_n263), .B(new_n303), .C1(new_n970), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n304), .A2(new_n286), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n851), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n951), .A2(new_n954), .A3(new_n836), .A4(new_n955), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n686), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  NOR4_X1   g791(.A1(new_n973), .A2(new_n975), .A3(new_n891), .A4(new_n977), .ZN(G57));
endmodule


