

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579;

  XNOR2_X1 U321 ( .A(n419), .B(n290), .ZN(n424) );
  INV_X1 U322 ( .A(n556), .ZN(n557) );
  NOR2_X1 U323 ( .A1(n488), .A2(n499), .ZN(n445) );
  AND2_X1 U324 ( .A1(G226GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U325 ( .A(n418), .B(n417), .Z(n290) );
  NOR2_X1 U326 ( .A1(n551), .A2(n453), .ZN(n454) );
  XNOR2_X1 U327 ( .A(G211GAT), .B(G218GAT), .ZN(n330) );
  NOR2_X1 U328 ( .A1(n509), .A2(n383), .ZN(n384) );
  XNOR2_X1 U329 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n462) );
  XNOR2_X1 U330 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U331 ( .A(n417), .B(n289), .ZN(n336) );
  XNOR2_X1 U332 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U333 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U334 ( .A(n569), .B(KEYINPUT41), .ZN(n556) );
  XNOR2_X1 U335 ( .A(n337), .B(n336), .ZN(n342) );
  INV_X1 U336 ( .A(G190GAT), .ZN(n470) );
  XNOR2_X1 U337 ( .A(n470), .B(KEYINPUT58), .ZN(n471) );
  XNOR2_X1 U338 ( .A(n446), .B(G99GAT), .ZN(n447) );
  XNOR2_X1 U339 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n448), .B(n447), .ZN(G1338GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n292) );
  XNOR2_X1 U342 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n306) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .Z(n334) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT77), .Z(n320) );
  XOR2_X1 U346 ( .A(n334), .B(n320), .Z(n294) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n295), .B(KEYINPUT72), .ZN(n420) );
  XOR2_X1 U351 ( .A(n420), .B(KEYINPUT11), .Z(n297) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT7), .B(KEYINPUT68), .Z(n301) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G29GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(KEYINPUT8), .B(n302), .Z(n444) );
  XOR2_X1 U359 ( .A(G50GAT), .B(G162GAT), .Z(n361) );
  XNOR2_X1 U360 ( .A(n444), .B(n361), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n551) );
  INV_X1 U363 ( .A(n551), .ZN(n469) );
  XNOR2_X1 U364 ( .A(KEYINPUT36), .B(n469), .ZN(n576) );
  XOR2_X1 U365 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n308) );
  XNOR2_X1 U366 ( .A(G127GAT), .B(KEYINPUT6), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U368 ( .A(KEYINPUT93), .B(KEYINPUT90), .Z(n310) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U371 ( .A(n312), .B(n311), .Z(n317) );
  XOR2_X1 U372 ( .A(KEYINPUT5), .B(G57GAT), .Z(n314) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT4), .B(n315), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n325) );
  XOR2_X1 U377 ( .A(G85GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(G120GAT), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n321) );
  XOR2_X1 U380 ( .A(n321), .B(n320), .Z(n323) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(G162GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U383 ( .A(n325), .B(n324), .Z(n329) );
  XNOR2_X1 U384 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n326), .B(KEYINPUT81), .ZN(n345) );
  XNOR2_X1 U386 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n327), .B(KEYINPUT2), .ZN(n368) );
  XNOR2_X1 U388 ( .A(n345), .B(n368), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n509) );
  XNOR2_X1 U390 ( .A(n330), .B(KEYINPUT21), .ZN(n331) );
  XOR2_X1 U391 ( .A(n331), .B(KEYINPUT87), .Z(n333) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n372) );
  XOR2_X1 U394 ( .A(n334), .B(n372), .Z(n337) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n335), .B(G64GAT), .ZN(n417) );
  XOR2_X1 U397 ( .A(G169GAT), .B(G8GAT), .Z(n432) );
  XOR2_X1 U398 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n339) );
  XNOR2_X1 U399 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(KEYINPUT19), .B(n340), .Z(n349) );
  XNOR2_X1 U402 ( .A(n432), .B(n349), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n511) );
  XOR2_X1 U404 ( .A(G176GAT), .B(KEYINPUT85), .Z(n344) );
  XNOR2_X1 U405 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n358) );
  XOR2_X1 U407 ( .A(G120GAT), .B(G71GAT), .Z(n414) );
  XOR2_X1 U408 ( .A(n414), .B(n345), .Z(n347) );
  NAND2_X1 U409 ( .A1(G227GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n356) );
  XOR2_X1 U412 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n351) );
  XNOR2_X1 U413 ( .A(G99GAT), .B(G134GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(n352), .B(G190GAT), .Z(n354) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G127GAT), .Z(n395) );
  XNOR2_X1 U417 ( .A(G43GAT), .B(n395), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n521) );
  NAND2_X1 U421 ( .A1(n511), .A2(n521), .ZN(n375) );
  XOR2_X1 U422 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n360) );
  XNOR2_X1 U423 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n365) );
  XOR2_X1 U425 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n363) );
  XOR2_X1 U426 ( .A(G141GAT), .B(G22GAT), .Z(n430) );
  XNOR2_X1 U427 ( .A(n430), .B(n361), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U429 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U430 ( .A1(G228GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U432 ( .A(n369), .B(n368), .Z(n374) );
  XOR2_X1 U433 ( .A(G78GAT), .B(G148GAT), .Z(n371) );
  XNOR2_X1 U434 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n418) );
  XNOR2_X1 U436 ( .A(n372), .B(n418), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n465) );
  NAND2_X1 U438 ( .A1(n375), .A2(n465), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n376), .B(KEYINPUT95), .ZN(n378) );
  XOR2_X1 U440 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n511), .B(KEYINPUT27), .ZN(n385) );
  NOR2_X1 U443 ( .A1(n465), .A2(n521), .ZN(n379) );
  XNOR2_X1 U444 ( .A(KEYINPUT26), .B(n379), .ZN(n563) );
  AND2_X1 U445 ( .A1(n385), .A2(n563), .ZN(n380) );
  NOR2_X1 U446 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n382), .B(KEYINPUT96), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(KEYINPUT97), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n509), .A2(n385), .ZN(n519) );
  NOR2_X1 U450 ( .A1(n521), .A2(n519), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n465), .B(KEYINPUT28), .ZN(n484) );
  NAND2_X1 U452 ( .A1(n386), .A2(n484), .ZN(n387) );
  NAND2_X1 U453 ( .A1(n388), .A2(n387), .ZN(n474) );
  XOR2_X1 U454 ( .A(G155GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U455 ( .A(G183GAT), .B(G71GAT), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U457 ( .A(n391), .B(G211GAT), .Z(n393) );
  XOR2_X1 U458 ( .A(G1GAT), .B(KEYINPUT69), .Z(n431) );
  XNOR2_X1 U459 ( .A(G22GAT), .B(n431), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n399) );
  XNOR2_X1 U461 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n394), .B(KEYINPUT70), .ZN(n413) );
  XOR2_X1 U463 ( .A(n413), .B(n395), .Z(n397) );
  NAND2_X1 U464 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(n399), .B(n398), .Z(n407) );
  XOR2_X1 U467 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n401) );
  XNOR2_X1 U468 ( .A(G8GAT), .B(G64GAT), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U470 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n403) );
  XNOR2_X1 U471 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n572) );
  NAND2_X1 U475 ( .A1(n474), .A2(n572), .ZN(n408) );
  NOR2_X1 U476 ( .A1(n576), .A2(n408), .ZN(n410) );
  XNOR2_X1 U477 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n410), .B(n409), .ZN(n488) );
  XOR2_X1 U479 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n412) );
  XNOR2_X1 U480 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n426) );
  XOR2_X1 U482 ( .A(KEYINPUT32), .B(n413), .Z(n416) );
  XNOR2_X1 U483 ( .A(n414), .B(G204GAT), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n419) );
  XOR2_X1 U485 ( .A(n420), .B(KEYINPUT75), .Z(n422) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n569) );
  XOR2_X1 U489 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n428) );
  NAND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n442) );
  XOR2_X1 U493 ( .A(G113GAT), .B(G197GAT), .Z(n434) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U496 ( .A(n435), .B(G36GAT), .Z(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n437) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(KEYINPUT30), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n438), .B(G50GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n565) );
  NAND2_X1 U504 ( .A1(n556), .A2(n565), .ZN(n499) );
  XOR2_X1 U505 ( .A(KEYINPUT105), .B(n445), .Z(n513) );
  NAND2_X1 U506 ( .A1(n513), .A2(n521), .ZN(n448) );
  XOR2_X1 U507 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n446) );
  INV_X1 U508 ( .A(n565), .ZN(n541) );
  NAND2_X1 U509 ( .A1(n556), .A2(n541), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n449) );
  XNOR2_X1 U511 ( .A(KEYINPUT110), .B(n449), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U513 ( .A1(n452), .A2(n572), .ZN(n453) );
  XNOR2_X1 U514 ( .A(KEYINPUT47), .B(n454), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n572), .A2(n576), .ZN(n456) );
  XNOR2_X1 U516 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n456), .B(n455), .ZN(n458) );
  AND2_X1 U518 ( .A1(n565), .A2(n569), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT48), .B(n461), .ZN(n518) );
  NAND2_X1 U522 ( .A1(n518), .A2(n511), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n509), .A2(n464), .ZN(n564) );
  NAND2_X1 U524 ( .A1(n564), .A2(n465), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT123), .B(KEYINPUT55), .Z(n466) );
  NAND2_X1 U526 ( .A1(n468), .A2(n521), .ZN(n560) );
  NOR2_X1 U527 ( .A1(n469), .A2(n560), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n541), .A2(n569), .ZN(n487) );
  NOR2_X1 U529 ( .A1(n572), .A2(n551), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT16), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n498) );
  NOR2_X1 U532 ( .A1(n487), .A2(n498), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(n476), .ZN(n485) );
  NAND2_X1 U534 ( .A1(n485), .A2(n509), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  XOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT99), .Z(n480) );
  NAND2_X1 U538 ( .A1(n511), .A2(n485), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n482) );
  NAND2_X1 U541 ( .A1(n485), .A2(n521), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n483), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n484), .ZN(n523) );
  NAND2_X1 U545 ( .A1(n485), .A2(n523), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U547 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U549 ( .A1(n496), .A2(n509), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n496), .A2(n511), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n496), .A2(n521), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U558 ( .A1(n523), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n501) );
  NOR2_X1 U561 ( .A1(n499), .A2(n498), .ZN(n506) );
  NAND2_X1 U562 ( .A1(n506), .A2(n509), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n506), .A2(n511), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n521), .A2(n506), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U571 ( .A1(n506), .A2(n523), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n513), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G92GAT), .ZN(G1337GAT) );
  XNOR2_X1 U577 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n517) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n523), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1339GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n525) );
  INV_X1 U583 ( .A(n518), .ZN(n520) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n539) );
  NAND2_X1 U585 ( .A1(n539), .A2(n521), .ZN(n522) );
  NOR2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n535), .A2(n541), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n528) );
  NAND2_X1 U591 ( .A1(n535), .A2(n556), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n531) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT115), .B(n532), .Z(n534) );
  INV_X1 U598 ( .A(n572), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n535), .A2(n547), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U602 ( .A1(n535), .A2(n551), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n539), .A2(n563), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT119), .B(n540), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n550), .A2(n541), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  NAND2_X1 U611 ( .A1(n550), .A2(n556), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT121), .Z(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n565), .A2(n560), .ZN(n553) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n553), .Z(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n560), .A2(n557), .ZN(n558) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(G1349GAT) );
  NOR2_X1 U626 ( .A1(n572), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n575) );
  NOR2_X1 U630 ( .A1(n565), .A2(n575), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n575), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n575), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(n573), .Z(n574) );
  XNOR2_X1 U639 ( .A(G211GAT), .B(n574), .ZN(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

