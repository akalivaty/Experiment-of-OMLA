//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT68), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G101), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n465), .B2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT3), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n471), .A2(G137), .A3(new_n462), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT69), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G137), .A4(new_n462), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n466), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(G160));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n473), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n462), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  NOR3_X1   g062(.A1(new_n481), .A2(new_n487), .A3(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT71), .B1(new_n476), .B2(new_n462), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(G136), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n471), .A2(new_n473), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n494), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n464), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n473), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n501), .B1(new_n506), .B2(new_n508), .ZN(G164));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(KEYINPUT77), .B1(G75), .B2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n515), .B1(KEYINPUT77), .B2(new_n514), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT75), .B(G651), .Z(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n512), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT76), .B(G88), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n519), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n519), .A2(new_n532), .A3(new_n526), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n527), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n525), .A2(G51), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n513), .A2(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n527), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n525), .A2(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n512), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n525), .A2(G43), .B1(new_n518), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n527), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT79), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n512), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n527), .A2(G91), .B1(G651), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n525), .A2(new_n567), .A3(G53), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n567), .B1(new_n525), .B2(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(G299));
  XNOR2_X1  g146(.A(new_n548), .B(KEYINPUT80), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  OR2_X1    g149(.A1(new_n513), .A2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n527), .A2(G87), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n525), .A2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G288));
  AND2_X1   g153(.A1(new_n513), .A2(G61), .ZN(new_n579));
  AND2_X1   g154(.A1(G73), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n518), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n521), .A2(new_n522), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(G48), .A3(G543), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n527), .A2(G86), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n527), .A2(KEYINPUT82), .A3(G86), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n585), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(G47), .A2(new_n525), .B1(new_n527), .B2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n512), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(new_n518), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n592), .A2(new_n599), .ZN(G290));
  XNOR2_X1  g175(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n583), .A2(new_n513), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n512), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n525), .A2(G54), .B1(G651), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  OR3_X1    g184(.A1(new_n602), .A2(new_n603), .A3(new_n601), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n572), .ZN(G284));
  AOI21_X1  g188(.A(new_n612), .B1(G868), .B2(new_n572), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n565), .A2(G651), .ZN(new_n616));
  INV_X1    g191(.A(G91), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n602), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n570), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n568), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n615), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(new_n611), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g204(.A1(new_n460), .A2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n464), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n490), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n482), .A2(G123), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(KEYINPUT85), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G111), .B2(new_n462), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n635), .B(new_n636), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n634), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT87), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n658), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  INV_X1    g243(.A(new_n665), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n669), .B2(new_n663), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n663), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n670), .B1(new_n673), .B2(new_n669), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n669), .A3(new_n666), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n683), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G16), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(G6), .A2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(G305), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G288), .B2(new_n701), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n702), .A2(new_n703), .ZN(new_n710));
  AND4_X1   g285(.A1(new_n699), .A2(new_n704), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n701), .A2(G24), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G290), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1986), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  OR2_X1    g293(.A1(G25), .A2(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n490), .A2(G131), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n482), .A2(G119), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n462), .A2(G107), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n719), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  AOI211_X1 g302(.A(new_n717), .B(new_n718), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n713), .B(new_n728), .C1(new_n726), .C2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n711), .A2(new_n712), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n729), .A2(KEYINPUT36), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT36), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n735), .B(new_n736), .Z(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  INV_X1    g313(.A(new_n464), .ZN(new_n739));
  INV_X1    g314(.A(G127), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n737), .B1(G2105), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n490), .A2(G139), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n725), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n725), .B2(G33), .ZN(new_n747));
  INV_X1    g322(.A(G2072), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n725), .A2(G32), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT26), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n630), .A2(G105), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n752), .B(new_n753), .C1(G129), .C2(new_n482), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n490), .A2(G141), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n747), .A2(new_n748), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n749), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n701), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n701), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G21), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G168), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n701), .A2(G19), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT91), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n555), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1341), .ZN(new_n775));
  INV_X1    g350(.A(G28), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n776), .B2(KEYINPUT30), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(KEYINPUT30), .B2(new_n776), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT31), .B(G11), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT95), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n778), .B(new_n780), .C1(new_n641), .C2(new_n725), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n764), .B2(new_n765), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n771), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n725), .A2(G27), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  INV_X1    g360(.A(new_n501), .ZN(new_n786));
  INV_X1    g361(.A(new_n508), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n507), .B1(new_n502), .B2(new_n504), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n785), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n762), .A2(new_n783), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G29), .A2(G35), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G162), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT29), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G2090), .Z(new_n797));
  NOR2_X1   g372(.A1(G4), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n623), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1348), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n725), .B1(new_n801), .B2(G34), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n801), .B2(G34), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G160), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2084), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n701), .A2(G20), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT23), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n725), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n490), .A2(G140), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n462), .A2(G116), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n482), .A2(G128), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(G29), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n800), .A2(new_n805), .A3(new_n810), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n793), .A2(new_n797), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n733), .A2(new_n824), .ZN(G311));
  INV_X1    g400(.A(G311), .ZN(G150));
  NAND2_X1  g401(.A1(new_n527), .A2(G93), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n525), .A2(G55), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n828), .C1(new_n517), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NOR2_X1   g407(.A1(new_n611), .A2(new_n624), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n555), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n832), .B1(new_n839), .B2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n756), .B(new_n819), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n724), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n482), .A2(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n462), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G142), .B2(new_n490), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n632), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n501), .A2(new_n505), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n744), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n745), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G160), .B(new_n641), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n857), .A2(new_n859), .A3(new_n862), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g443(.A(G166), .B(G305), .Z(new_n869));
  XNOR2_X1  g444(.A(G290), .B(G288), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  OR3_X1    g448(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n626), .B(new_n836), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n611), .B(G299), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n611), .B(new_n620), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n892), .B2(new_n889), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n885), .B1(new_n893), .B2(new_n883), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n882), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n880), .A2(new_n894), .A3(new_n881), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  MUX2_X1   g473(.A(new_n830), .B(new_n898), .S(G868), .Z(G295));
  MUX2_X1   g474(.A(new_n830), .B(new_n898), .S(G868), .Z(G331));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND3_X1  g476(.A1(G171), .A2(KEYINPUT102), .A3(G286), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(G168), .B2(new_n548), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n902), .B(new_n904), .C1(new_n572), .C2(G286), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(new_n836), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n893), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n884), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n876), .ZN(new_n911));
  INV_X1    g486(.A(new_n876), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n901), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n892), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n915), .A2(new_n906), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n876), .B1(new_n916), .B2(new_n908), .ZN(new_n917));
  AND4_X1   g492(.A1(new_n901), .A2(new_n913), .A3(new_n865), .A4(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n914), .A2(new_n918), .A3(KEYINPUT44), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n901), .A3(new_n913), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n913), .A2(new_n865), .A3(new_n917), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n901), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(KEYINPUT44), .B2(new_n922), .ZN(G397));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n501), .B2(new_n505), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n478), .A2(new_n475), .ZN(new_n928));
  NAND2_X1  g503(.A1(G113), .A2(G2104), .ZN(new_n929));
  INV_X1    g504(.A(G125), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n739), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n931), .A2(G2105), .B1(G101), .B2(new_n630), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n928), .A2(new_n932), .A3(G40), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n756), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n819), .B(new_n821), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT104), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n724), .B(new_n727), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n934), .A2(G290), .A3(G1986), .ZN(new_n945));
  INV_X1    g520(.A(new_n934), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n716), .B1(new_n592), .B2(new_n599), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT103), .Z(new_n949));
  AND2_X1   g524(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT54), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT45), .B1(new_n789), .B2(new_n924), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT45), .B(new_n924), .C1(new_n501), .C2(new_n505), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n933), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n791), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n479), .A2(G40), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n926), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n958), .A2(new_n959), .B1(new_n765), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n927), .A2(new_n960), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n789), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n971), .A2(new_n572), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n968), .A2(KEYINPUT53), .A3(new_n791), .A4(new_n953), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n572), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n951), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G2084), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n964), .A2(new_n977), .B1(new_n970), .B2(new_n766), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G286), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n978), .B2(G168), .ZN(new_n983));
  NAND2_X1  g558(.A1(KEYINPUT127), .A2(KEYINPUT51), .ZN(new_n984));
  OR2_X1    g559(.A1(KEYINPUT127), .A2(KEYINPUT51), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n984), .B2(new_n983), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n974), .A2(G171), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(KEYINPUT54), .C1(new_n572), .C2(new_n971), .ZN(new_n990));
  NAND2_X1  g565(.A1(G303), .A2(G8), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT107), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR4_X1    g568(.A1(KEYINPUT107), .A2(G166), .A3(new_n992), .A4(new_n979), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n955), .B(KEYINPUT106), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n698), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n925), .A2(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n933), .A2(new_n999), .A3(KEYINPUT114), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n789), .A2(new_n961), .A3(new_n924), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT114), .B1(new_n933), .B2(new_n999), .ZN(new_n1003));
  OR3_X1    g578(.A1(new_n1002), .A2(G2090), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n979), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n996), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(G8), .B1(new_n960), .B2(new_n925), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1008), .B(new_n1009), .C1(new_n1010), .C2(G288), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT108), .B(G1976), .ZN(new_n1012));
  AND2_X1   g587(.A1(G288), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(new_n1013), .B2(new_n1008), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1011), .B(new_n1014), .Z(new_n1015));
  NOR2_X1   g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n586), .A2(new_n581), .A3(new_n584), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(KEYINPUT110), .A3(G1981), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(G1981), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1019), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n1016), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1026), .A3(new_n1008), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT111), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1023), .A2(new_n1026), .A3(new_n1029), .A4(new_n1008), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1015), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n998), .B1(G2090), .B2(new_n965), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n996), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1006), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n976), .A2(new_n988), .A3(new_n990), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n623), .A2(KEYINPUT125), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n960), .A2(new_n925), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n821), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT119), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n964), .A2(G1348), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n611), .B(KEYINPUT125), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(KEYINPUT60), .A3(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1045), .B(new_n1047), .C1(KEYINPUT60), .C2(new_n1042), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n809), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(G164), .B2(G1384), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n933), .A3(new_n953), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n954), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(KEYINPUT118), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT115), .B(new_n809), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1052), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(KEYINPUT57), .C1(new_n620), .C2(KEYINPUT116), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(G299), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(new_n1052), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT123), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1079), .A3(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1072), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n952), .A2(new_n954), .A3(G1996), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT58), .B(G1341), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1083), .A2(KEYINPUT121), .B1(new_n1038), .B2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n955), .A2(KEYINPUT121), .A3(new_n935), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n556), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT59), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(new_n556), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1082), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1049), .B1(new_n1081), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1079), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT123), .B(new_n1075), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1092), .B(new_n1049), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1048), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1073), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1043), .A2(new_n623), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1072), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n1101), .B(KEYINPUT120), .Z(new_n1102));
  AOI21_X1  g677(.A(new_n1036), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n982), .A2(new_n987), .A3(KEYINPUT62), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT62), .B1(new_n982), .B2(new_n987), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(new_n972), .A3(new_n1035), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT63), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n980), .A2(G168), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1034), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1107), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1032), .A2(G8), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n996), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1031), .A2(new_n1112), .A3(new_n996), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT112), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1017), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1007), .B1(new_n1120), .B2(KEYINPUT113), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1122), .A3(new_n1017), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1106), .A2(new_n1114), .A3(new_n1115), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n950), .B1(new_n1103), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n937), .A2(new_n755), .A3(new_n754), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n934), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT46), .B1(new_n934), .B2(G1996), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1127), .A2(new_n946), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT47), .ZN(new_n1131));
  INV_X1    g706(.A(new_n727), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n724), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n939), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n814), .A2(new_n821), .A3(new_n818), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n934), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n945), .B(KEYINPUT48), .Z(new_n1137));
  AOI211_X1 g712(.A(new_n1131), .B(new_n1136), .C1(new_n944), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1126), .A2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g714(.A1(new_n914), .A2(new_n918), .ZN(new_n1141));
  INV_X1    g715(.A(G319), .ZN(new_n1142));
  NOR4_X1   g716(.A1(G401), .A2(new_n1142), .A3(G227), .A4(G229), .ZN(new_n1143));
  AND3_X1   g717(.A1(new_n1141), .A2(new_n867), .A3(new_n1143), .ZN(G308));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n867), .A3(new_n1143), .ZN(G225));
endmodule


