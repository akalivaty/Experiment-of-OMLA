//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n193), .B2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT23), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n192), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(new_n194), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n203), .B2(G110), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT80), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(KEYINPUT78), .A3(G140), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(KEYINPUT78), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT79), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n212));
  INV_X1    g026(.A(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n217), .B2(new_n212), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT16), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n213), .A3(G125), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n211), .A2(new_n220), .A3(G146), .A4(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n205), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n221), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n219), .B1(new_n218), .B2(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n222), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n195), .A2(new_n196), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n203), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n203), .A2(new_n232), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(G110), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n225), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT22), .B(G137), .ZN(new_n239));
  INV_X1    g053(.A(G953), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n240), .A2(G221), .A3(G234), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n239), .B(new_n241), .Z(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n225), .B(new_n242), .C1(new_n231), .C2(new_n237), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n188), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT81), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n244), .A2(new_n188), .A3(new_n245), .A4(new_n248), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n190), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n244), .A2(new_n245), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n253), .A2(G902), .A3(new_n189), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G237), .ZN(new_n260));
  AOI21_X1  g074(.A(G953), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n223), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G146), .ZN(new_n272));
  AND4_X1   g086(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(G146), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n223), .B2(G143), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(KEYINPUT64), .A3(G146), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n191), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n279));
  OAI22_X1  g093(.A1(new_n269), .A2(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G134), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G137), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT11), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n284), .B2(G137), .ZN(new_n290));
  AOI21_X1  g104(.A(G131), .B1(new_n284), .B2(G137), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n282), .A2(KEYINPUT11), .A3(G134), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT69), .B1(new_n295), .B2(new_n286), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n280), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G116), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n193), .A2(G116), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G113), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n303), .A2(new_n304), .A3(new_n310), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n290), .A2(new_n292), .A3(new_n285), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G131), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n293), .ZN(new_n317));
  AND2_X1   g131(.A1(KEYINPUT0), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n267), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT0), .A2(G128), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n278), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n314), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n280), .A2(new_n325), .A3(new_n294), .A4(new_n296), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n298), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT71), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n298), .A2(new_n329), .A3(new_n324), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n287), .A2(new_n293), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n267), .A2(new_n266), .A3(new_n268), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n271), .A2(KEYINPUT64), .A3(G146), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT64), .B1(new_n271), .B2(G146), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n270), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n279), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n332), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(KEYINPUT65), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT65), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n344), .B(new_n319), .C1(new_n278), .C2(new_n321), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n317), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n342), .B1(new_n346), .B2(KEYINPUT66), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n343), .A2(new_n348), .A3(new_n317), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n314), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n331), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT28), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n324), .A2(new_n297), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n265), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n331), .A2(KEYINPUT73), .A3(new_n265), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT30), .B1(new_n347), .B2(new_n349), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n323), .A2(new_n317), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n298), .A2(KEYINPUT30), .A3(new_n362), .A4(new_n326), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n314), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT31), .ZN(new_n366));
  INV_X1    g180(.A(new_n265), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n328), .B2(new_n330), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n363), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n360), .ZN(new_n372));
  AOI22_X1  g186(.A1(KEYINPUT73), .A2(new_n368), .B1(new_n372), .B2(new_n314), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n331), .A2(new_n265), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT31), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n358), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n379));
  NOR2_X1   g193(.A1(G472), .A2(G902), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n366), .B1(new_n365), .B2(new_n369), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(KEYINPUT31), .A3(new_n364), .A4(new_n359), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n357), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n380), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT32), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n367), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n298), .A2(new_n362), .A3(new_n326), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n328), .A2(new_n330), .B1(new_n314), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n356), .B(new_n390), .C1(new_n392), .C2(new_n355), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n188), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n328), .A2(new_n330), .B1(new_n350), .B2(new_n314), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n356), .B(new_n265), .C1(new_n395), .C2(new_n355), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n364), .A2(new_n331), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n397), .B2(new_n367), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G472), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n388), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n393), .A2(new_n188), .ZN(new_n402));
  INV_X1    g216(.A(new_n314), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n371), .A2(new_n360), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n331), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n367), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n396), .A3(new_n389), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n400), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n256), .B1(new_n387), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n304), .A2(KEYINPUT5), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n306), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n305), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G104), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(new_n416), .B2(G107), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G104), .ZN(new_n420));
  INV_X1    g234(.A(G101), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(G107), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n419), .A2(G104), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n416), .A2(G107), .ZN(new_n425));
  OAI21_X1  g239(.A(G101), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n415), .A2(new_n313), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G101), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT4), .A3(new_n423), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(G101), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n303), .A2(new_n304), .A3(new_n310), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n310), .B1(new_n303), .B2(new_n304), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n428), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT90), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n314), .A2(new_n431), .A3(new_n434), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n428), .ZN(new_n442));
  XOR2_X1   g256(.A(G110), .B(G122), .Z(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n428), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(KEYINPUT6), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n322), .A2(G125), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT91), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n336), .A2(new_n341), .A3(new_n206), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n322), .A2(new_n452), .A3(G125), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G224), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G953), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n439), .A2(new_n458), .A3(new_n442), .A4(new_n443), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n443), .B(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n428), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n427), .B1(new_n415), .B2(new_n313), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n451), .A2(new_n449), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n456), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n456), .A2(new_n467), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n450), .A2(new_n451), .A3(new_n453), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n465), .A2(new_n468), .A3(new_n470), .A4(new_n446), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n471), .A2(new_n188), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n460), .A2(new_n472), .A3(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G214), .B1(G237), .B2(G902), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n240), .A2(G952), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT99), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n478), .A2(new_n479), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G478), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT9), .B(G234), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n493), .A2(new_n187), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n271), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n191), .A2(G143), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n284), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n271), .A2(KEYINPUT13), .A3(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n497), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n191), .B2(G143), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT97), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n496), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n498), .B1(new_n506), .B2(new_n284), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n300), .A2(new_n302), .A3(G122), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n299), .A2(G122), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n419), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT96), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(G107), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n507), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G107), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n496), .A2(new_n497), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G134), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n498), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n508), .A2(new_n523), .A3(new_n510), .ZN(new_n524));
  OAI21_X1  g338(.A(G107), .B1(new_n508), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n495), .B1(new_n518), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n507), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n511), .A2(new_n512), .A3(new_n419), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(new_n519), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n513), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n494), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT98), .B1(new_n534), .B2(new_n188), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT98), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n536), .B(G902), .C1(new_n528), .C2(new_n533), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n492), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n188), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n491), .B(G478), .C1(new_n539), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G475), .A2(G902), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n259), .A2(G237), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n545));
  OAI211_X1 g359(.A(G214), .B(new_n240), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n271), .ZN(new_n547));
  AOI21_X1  g361(.A(G143), .B1(new_n261), .B2(G214), .ZN(new_n548));
  OAI21_X1  g362(.A(G131), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n271), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n281), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n281), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n228), .A2(new_n554), .A3(new_n222), .A4(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT18), .B(G131), .C1(new_n547), .C2(new_n548), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n224), .B1(new_n218), .B2(new_n223), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT18), .A2(G131), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n551), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G113), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n416), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n557), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n551), .A2(new_n281), .A3(new_n552), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT93), .B1(new_n566), .B2(new_n555), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n549), .A2(new_n568), .A3(new_n553), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n217), .A2(new_n570), .A3(KEYINPUT95), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n209), .A2(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT95), .B1(new_n217), .B2(new_n570), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n571), .A2(new_n572), .A3(new_n223), .A4(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n567), .A2(new_n222), .A3(new_n569), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n564), .B1(new_n575), .B2(new_n562), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n543), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT20), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n579), .B(new_n543), .C1(new_n565), .C2(new_n576), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n564), .B1(new_n557), .B2(new_n562), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n188), .B1(new_n565), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n578), .A2(new_n580), .B1(G475), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n542), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n490), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G221), .ZN(new_n586));
  INV_X1    g400(.A(new_n493), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n188), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n240), .A2(G227), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT82), .ZN(new_n591));
  XNOR2_X1  g405(.A(G110), .B(G140), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n267), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT84), .B(KEYINPUT1), .C1(new_n271), .C2(G146), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G128), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT84), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT85), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(new_n594), .C1(new_n596), .C2(new_n597), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n336), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT10), .B1(new_n602), .B2(new_n427), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n427), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n323), .A2(new_n431), .A3(new_n434), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n317), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n593), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT86), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT12), .B1(new_n317), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n423), .A2(new_n426), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n336), .A2(new_n341), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n602), .B2(new_n427), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(new_n608), .ZN(new_n615));
  INV_X1    g429(.A(new_n611), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n598), .A2(KEYINPUT85), .B1(new_n335), .B2(new_n334), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n612), .B1(new_n617), .B2(new_n601), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n317), .B(new_n616), .C1(new_n618), .C2(new_n613), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n602), .A2(new_n427), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n606), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n608), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n603), .A2(new_n606), .A3(new_n317), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n593), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT88), .B(G469), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n629), .A2(KEYINPUT89), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT89), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G469), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n593), .B(KEYINPUT83), .Z(new_n635));
  INV_X1    g449(.A(new_n627), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n635), .B1(new_n620), .B2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n626), .A2(new_n627), .A3(new_n593), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT87), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n317), .B1(new_n603), .B2(new_n606), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n609), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT87), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n627), .B1(new_n619), .B2(new_n615), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n635), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n634), .B1(new_n645), .B2(new_n188), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n589), .B1(new_n633), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n585), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n411), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G101), .ZN(G3));
  OAI21_X1  g464(.A(G472), .B1(new_n384), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n378), .A2(new_n380), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n647), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n539), .A2(G478), .ZN(new_n655));
  AND2_X1   g469(.A1(G478), .A2(G902), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n534), .A2(KEYINPUT33), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n534), .A2(KEYINPUT33), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(G478), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n583), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n476), .A2(new_n664), .A3(new_n477), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n460), .A2(KEYINPUT100), .A3(new_n472), .A4(new_n474), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n479), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n663), .A2(new_n488), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n654), .A2(new_n255), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT34), .B(G104), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n578), .A2(new_n673), .A3(new_n580), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n582), .A2(G475), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n577), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n541), .A4(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n668), .A2(new_n677), .A3(new_n488), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n654), .A2(new_n255), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT102), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT103), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  XNOR2_X1  g497(.A(new_n238), .B(KEYINPUT104), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n243), .A2(KEYINPUT36), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n238), .A2(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n238), .A2(KEYINPUT104), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n189), .A2(G902), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n252), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n585), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n654), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT37), .B(G110), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT105), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n695), .B(new_n697), .ZN(G12));
  AOI21_X1  g512(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n384), .A2(KEYINPUT32), .A3(new_n385), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n388), .B(new_n400), .C1(new_n402), .C2(new_n407), .ZN(new_n702));
  OAI22_X1  g516(.A1(new_n699), .A2(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n240), .A2(G900), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(G902), .A3(new_n481), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n483), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n668), .A2(new_n677), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n647), .B1(new_n709), .B2(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n250), .A2(new_n251), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n189), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n687), .A2(new_n690), .A3(new_n692), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n677), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n666), .A2(new_n479), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n460), .A2(new_n472), .A3(new_n474), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n474), .B1(new_n460), .B2(new_n472), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n716), .B1(new_n719), .B2(new_n664), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n715), .A2(new_n720), .A3(new_n707), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n703), .A2(new_n710), .A3(new_n714), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  NAND2_X1  g539(.A1(new_n645), .A2(new_n188), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n621), .A2(new_n628), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n188), .A3(new_n630), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n629), .A2(KEYINPUT89), .A3(new_n630), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n588), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n707), .B(KEYINPUT39), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n392), .A2(new_n265), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n373), .B2(new_n376), .ZN(new_n740));
  OAI21_X1  g554(.A(G472), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n387), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n478), .B(KEYINPUT38), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n542), .A2(new_n583), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n479), .A2(new_n693), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n737), .A2(new_n738), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G143), .ZN(G45));
  NAND4_X1  g561(.A1(new_n720), .A2(KEYINPUT108), .A3(new_n662), .A4(new_n707), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n578), .A2(new_n580), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n675), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n657), .A2(new_n660), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n707), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n749), .B1(new_n753), .B2(new_n668), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n703), .A2(new_n734), .A3(new_n714), .A4(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT109), .B(G146), .Z(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G48));
  OR2_X1    g572(.A1(new_n629), .A2(new_n634), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n589), .B(new_n759), .C1(new_n631), .C2(new_n632), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT110), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n703), .A2(new_n761), .A3(new_n255), .A4(new_n669), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT41), .B(G113), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NAND4_X1  g578(.A1(new_n703), .A2(new_n761), .A3(new_n255), .A4(new_n678), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G116), .ZN(G18));
  NOR4_X1   g580(.A1(new_n760), .A2(new_n668), .A3(new_n584), .A4(new_n488), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n703), .A2(new_n714), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  OAI21_X1  g583(.A(new_n356), .B1(new_n392), .B2(new_n355), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n367), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n370), .B2(new_n377), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n380), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n651), .A2(new_n773), .A3(new_n255), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n720), .A2(new_n744), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n488), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n761), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  NAND3_X1  g592(.A1(new_n651), .A2(new_n773), .A3(new_n714), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n760), .A2(new_n668), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n753), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n662), .A2(KEYINPUT111), .A3(new_n707), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  OAI21_X1  g602(.A(new_n641), .B1(new_n643), .B2(new_n635), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n188), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(G469), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n733), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n479), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n588), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n478), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n703), .A2(new_n255), .A3(new_n786), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(KEYINPUT112), .A2(KEYINPUT42), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n800), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n411), .A2(new_n786), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  NOR2_X1   g619(.A1(new_n677), .A2(new_n708), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n703), .A2(new_n255), .A3(new_n798), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n284), .ZN(G36));
  NAND2_X1  g622(.A1(G469), .A2(G902), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT45), .B1(new_n639), .B2(new_n644), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n789), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT46), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n633), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n816), .A2(new_n589), .A3(new_n735), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n478), .A2(new_n793), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT114), .Z(new_n819));
  NAND2_X1  g633(.A1(new_n752), .A2(new_n583), .ZN(new_n820));
  NOR2_X1   g634(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n820), .B1(new_n823), .B2(new_n821), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n653), .A2(new_n714), .A3(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT44), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT44), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n817), .B(new_n819), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(KEYINPUT115), .B(G137), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(G39));
  AND3_X1   g645(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n589), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT47), .B1(new_n816), .B2(new_n589), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n818), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n703), .A2(new_n255), .A3(new_n753), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  AOI21_X1  g652(.A(new_n483), .B1(new_n822), .B2(new_n824), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n774), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n743), .A2(new_n479), .A3(new_n760), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT50), .Z(new_n843));
  OR2_X1    g657(.A1(new_n835), .A2(new_n760), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n742), .A2(new_n256), .A3(new_n844), .A4(new_n483), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n583), .A2(new_n661), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n839), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n844), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n845), .A2(new_n847), .B1(new_n849), .B2(new_n780), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n733), .A2(new_n759), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n589), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT117), .B1(new_n834), .B2(new_n855), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n819), .A3(new_n840), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n853), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n840), .A2(new_n781), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n480), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n849), .A2(new_n411), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT48), .Z(new_n864));
  AOI211_X1 g678(.A(new_n862), .B(new_n864), .C1(new_n662), .C2(new_n845), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n853), .B(new_n866), .C1(new_n856), .C2(new_n858), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n840), .A2(new_n819), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n834), .A2(KEYINPUT116), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n855), .B1(new_n834), .B2(KEYINPUT116), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n852), .B1(new_n871), .B2(new_n851), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n860), .A2(new_n865), .A3(new_n867), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(new_n653), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n583), .A2(new_n541), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n490), .B1(new_n663), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n255), .A3(new_n734), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n768), .A2(new_n878), .A3(new_n777), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n779), .A2(new_n785), .A3(new_n797), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n647), .B(new_n693), .C1(new_n387), .C2(new_n410), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n542), .A2(new_n675), .A3(new_n707), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n674), .A2(new_n676), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n835), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n411), .A2(new_n648), .B1(new_n654), .B2(new_n694), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n411), .B(new_n761), .C1(new_n669), .C2(new_n678), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n879), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n807), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n804), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n712), .A2(new_n589), .A3(new_n713), .A4(new_n707), .ZN(new_n892));
  INV_X1    g706(.A(new_n792), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n775), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n742), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n724), .A2(new_n756), .A3(new_n787), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n715), .A2(new_n720), .A3(KEYINPUT107), .A4(new_n707), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n734), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n668), .A2(new_n677), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT107), .B1(new_n900), .B2(new_n707), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n693), .B1(new_n387), .B2(new_n410), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n779), .A2(new_n785), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(new_n781), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n756), .A4(new_n895), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n897), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n891), .B(new_n908), .C1(KEYINPUT53), .C2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n807), .B1(new_n801), .B2(new_n803), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n649), .A2(new_n762), .A3(new_n765), .A4(new_n695), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n879), .A4(new_n885), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n897), .A2(new_n907), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n874), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT53), .B1(new_n891), .B2(new_n908), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT53), .B1(new_n905), .B2(new_n906), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n914), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n873), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n255), .A2(new_n583), .A3(new_n752), .A4(new_n794), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT49), .ZN(new_n926));
  INV_X1    g740(.A(new_n854), .ZN(new_n927));
  AOI211_X1 g741(.A(new_n743), .B(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n923), .A2(new_n924), .B1(new_n742), .B2(new_n929), .ZN(G75));
  NOR2_X1   g744(.A1(new_n240), .A2(G952), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n919), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n891), .A2(new_n908), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n188), .B1(new_n934), .B2(new_n916), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(G210), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n448), .A2(new_n459), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n457), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n932), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n916), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(G902), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n475), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n941), .B1(new_n948), .B2(new_n950), .ZN(G51));
  XOR2_X1   g765(.A(new_n809), .B(KEYINPUT57), .Z(new_n952));
  AOI21_X1  g766(.A(new_n874), .B1(new_n934), .B2(new_n916), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n921), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT121), .B(new_n952), .C1(new_n921), .C2(new_n953), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n728), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n810), .A2(new_n812), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n947), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n931), .B1(new_n958), .B2(new_n960), .ZN(G54));
  AND2_X1   g775(.A1(KEYINPUT58), .A2(G475), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n945), .A2(new_n946), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n565), .A2(new_n576), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n931), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n945), .A2(new_n966), .A3(new_n946), .A4(new_n962), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(G60));
  NAND2_X1  g782(.A1(new_n658), .A2(new_n659), .ZN(new_n969));
  XOR2_X1   g783(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n656), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n922), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n969), .B(new_n971), .C1(new_n921), .C2(new_n953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n932), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT123), .B1(new_n942), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n980), .B(new_n977), .C1(new_n934), .C2(new_n916), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n691), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n918), .B2(new_n920), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n980), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n942), .A2(KEYINPUT123), .A3(new_n978), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n253), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n982), .A2(new_n986), .A3(new_n932), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n982), .A2(new_n986), .A3(KEYINPUT61), .A4(new_n932), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  OAI21_X1  g805(.A(G953), .B1(new_n485), .B2(new_n455), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n913), .A2(new_n879), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(G953), .ZN(new_n994));
  INV_X1    g808(.A(G898), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n937), .B1(new_n995), .B2(G953), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n994), .B(new_n996), .Z(G69));
  NAND3_X1  g811(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n372), .B(new_n998), .Z(new_n999));
  AOI21_X1  g813(.A(new_n835), .B1(new_n663), .B2(new_n876), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n411), .A2(new_n734), .A3(new_n735), .A4(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n837), .A2(new_n829), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n905), .A2(new_n756), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n746), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(new_n1006), .A3(new_n746), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1002), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n999), .B1(new_n1008), .B2(new_n240), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT124), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n1011), .B(new_n999), .C1(new_n1008), .C2(new_n240), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n817), .A2(new_n411), .A3(new_n720), .A4(new_n744), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n837), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1003), .A2(new_n829), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT125), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1003), .A2(new_n829), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1015), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n912), .B(KEYINPUT126), .ZN(new_n1021));
  AOI21_X1  g835(.A(G953), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n999), .B1(new_n1022), .B2(new_n704), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n240), .B1(G227), .B2(G900), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1013), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1013), .B2(new_n1023), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1025), .A2(new_n1026), .ZN(G72));
  OAI21_X1  g841(.A(new_n406), .B1(new_n365), .B2(new_n369), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(new_n910), .B2(new_n916), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT127), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1020), .A2(new_n993), .A3(new_n1021), .ZN(new_n1034));
  AOI211_X1 g848(.A(new_n265), .B(new_n397), .C1(new_n1034), .C2(new_n1030), .ZN(new_n1035));
  INV_X1    g849(.A(new_n993), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1030), .B1(new_n1008), .B2(new_n1036), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1037), .A2(new_n265), .A3(new_n397), .ZN(new_n1038));
  NOR4_X1   g852(.A1(new_n1033), .A2(new_n1035), .A3(new_n1038), .A4(new_n931), .ZN(G57));
endmodule


