

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G651), .A2(n594), .ZN(n804) );
  NAND2_X1 U555 ( .A1(n626), .A2(n625), .ZN(n789) );
  AND2_X2 U556 ( .A1(n639), .A2(G1341), .ZN(n627) );
  NOR2_X2 U557 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X2 U558 ( .A1(G543), .A2(n544), .ZN(n536) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n799) );
  NOR2_X4 U560 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  NOR2_X1 U561 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X2 U562 ( .A1(G2104), .A2(n527), .ZN(n888) );
  BUF_X1 U563 ( .A(n799), .Z(n523) );
  XNOR2_X1 U564 ( .A(n532), .B(KEYINPUT65), .ZN(n553) );
  INV_X1 U565 ( .A(KEYINPUT0), .ZN(n538) );
  NAND2_X1 U566 ( .A1(n553), .A2(G101), .ZN(n533) );
  XNOR2_X1 U567 ( .A(n552), .B(n551), .ZN(G168) );
  XNOR2_X1 U568 ( .A(KEYINPUT75), .B(KEYINPUT7), .ZN(n551) );
  OR2_X1 U569 ( .A1(n951), .A2(n645), .ZN(n524) );
  AND2_X1 U570 ( .A1(n724), .A2(G137), .ZN(n525) );
  INV_X1 U571 ( .A(KEYINPUT27), .ZN(n608) );
  XNOR2_X1 U572 ( .A(n609), .B(n608), .ZN(n611) );
  BUF_X1 U573 ( .A(n639), .Z(n671) );
  OR2_X1 U574 ( .A1(n670), .A2(n691), .ZN(n678) );
  AND2_X1 U575 ( .A1(n678), .A2(n677), .ZN(n679) );
  INV_X1 U576 ( .A(KEYINPUT32), .ZN(n681) );
  INV_X1 U577 ( .A(n965), .ZN(n699) );
  NOR2_X1 U578 ( .A1(n713), .A2(n699), .ZN(n700) );
  INV_X1 U579 ( .A(n953), .ZN(n705) );
  INV_X1 U580 ( .A(KEYINPUT97), .ZN(n717) );
  BUF_X1 U581 ( .A(n616), .Z(n803) );
  XNOR2_X1 U582 ( .A(KEYINPUT73), .B(KEYINPUT5), .ZN(n547) );
  XNOR2_X1 U583 ( .A(n538), .B(G543), .ZN(n594) );
  BUF_X1 U584 ( .A(n620), .Z(n800) );
  XNOR2_X1 U585 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U586 ( .A(KEYINPUT67), .B(n582), .Z(G171) );
  XOR2_X1 U587 ( .A(KEYINPUT17), .B(n526), .Z(n724) );
  INV_X1 U588 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U589 ( .A1(G125), .A2(n888), .ZN(n529) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U591 ( .A1(G113), .A2(n889), .ZN(n528) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n525), .A2(n530), .ZN(n535) );
  INV_X1 U594 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n531), .A2(G2104), .ZN(n532) );
  XOR2_X1 U596 ( .A(n533), .B(KEYINPUT23), .Z(n534) );
  AND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(G160) );
  INV_X1 U598 ( .A(G651), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n536), .Z(n620) );
  NAND2_X1 U600 ( .A1(n800), .A2(G63), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(KEYINPUT74), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G51), .A2(n804), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT6), .B(n541), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G89), .A2(n523), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT4), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(KEYINPUT72), .ZN(n546) );
  NOR2_X1 U608 ( .A1(n594), .A2(n544), .ZN(n616) );
  NAND2_X1 U609 ( .A1(G76), .A2(n803), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n552) );
  BUF_X2 U612 ( .A(n553), .Z(n723) );
  NAND2_X1 U613 ( .A1(G102), .A2(n723), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G138), .A2(n724), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G126), .A2(n888), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G114), .A2(n889), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X2 U619 ( .A1(n559), .A2(n558), .ZN(G164) );
  NAND2_X1 U620 ( .A1(G73), .A2(n803), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT2), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G61), .A2(n800), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G48), .A2(n804), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n523), .A2(G86), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT80), .B(n563), .Z(n564) );
  NOR2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(G305) );
  NAND2_X1 U629 ( .A1(G91), .A2(n523), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G78), .A2(n803), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n800), .A2(G65), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT68), .B(n570), .Z(n571) );
  NOR2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n804), .A2(G53), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(G299) );
  NAND2_X1 U637 ( .A1(G64), .A2(n800), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G52), .A2(n804), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G90), .A2(n523), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G77), .A2(n803), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n579), .Z(n580) );
  NOR2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U645 ( .A(G171), .ZN(G301) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT76), .B(n583), .ZN(G286) );
  NAND2_X1 U648 ( .A1(G88), .A2(n523), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G75), .A2(n803), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G50), .A2(n804), .ZN(n586) );
  XNOR2_X1 U652 ( .A(KEYINPUT81), .B(n586), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n800), .A2(G62), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(G303) );
  NAND2_X1 U656 ( .A1(G49), .A2(n804), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G74), .A2(G651), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U659 ( .A1(n800), .A2(n593), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n594), .A2(G87), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(G288) );
  NAND2_X1 U662 ( .A1(G85), .A2(n523), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G72), .A2(n803), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U665 ( .A1(G47), .A2(n804), .ZN(n599) );
  XOR2_X1 U666 ( .A(KEYINPUT66), .B(n599), .Z(n600) );
  NOR2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n800), .A2(G60), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(G290) );
  NAND2_X1 U670 ( .A1(G160), .A2(G40), .ZN(n721) );
  INV_X1 U671 ( .A(n721), .ZN(n604) );
  NOR2_X2 U672 ( .A1(G164), .A2(G1384), .ZN(n722) );
  NAND2_X2 U673 ( .A1(n604), .A2(n722), .ZN(n639) );
  NAND2_X1 U674 ( .A1(G8), .A2(n639), .ZN(n713) );
  NOR2_X1 U675 ( .A1(G1981), .A2(G305), .ZN(n605) );
  XOR2_X1 U676 ( .A(n605), .B(KEYINPUT24), .Z(n606) );
  NOR2_X1 U677 ( .A1(n713), .A2(n606), .ZN(n720) );
  INV_X1 U678 ( .A(n639), .ZN(n656) );
  INV_X1 U679 ( .A(KEYINPUT91), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n656), .B(n607), .ZN(n638) );
  NAND2_X1 U681 ( .A1(n638), .A2(G2072), .ZN(n609) );
  INV_X1 U682 ( .A(n638), .ZN(n655) );
  NAND2_X1 U683 ( .A1(G1956), .A2(n655), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n647) );
  NAND2_X1 U685 ( .A1(G299), .A2(n647), .ZN(n612) );
  XOR2_X1 U686 ( .A(KEYINPUT28), .B(n612), .Z(n653) );
  INV_X1 U687 ( .A(n639), .ZN(n613) );
  AND2_X1 U688 ( .A1(n613), .A2(G1996), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT26), .ZN(n629) );
  NAND2_X1 U690 ( .A1(n799), .A2(G81), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT12), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G68), .A2(n616), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT13), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n620), .A2(G56), .ZN(n621) );
  XNOR2_X1 U696 ( .A(KEYINPUT14), .B(n621), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(KEYINPUT71), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n804), .A2(G43), .ZN(n625) );
  OR2_X2 U700 ( .A1(n627), .A2(n789), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U702 ( .A1(G92), .A2(n523), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G66), .A2(n800), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U705 ( .A1(G79), .A2(n803), .ZN(n634) );
  NAND2_X1 U706 ( .A1(G54), .A2(n804), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U709 ( .A(KEYINPUT15), .B(n637), .Z(n951) );
  NAND2_X1 U710 ( .A1(n645), .A2(n951), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n638), .A2(G2067), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G1348), .A2(n671), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n644), .B(KEYINPUT92), .ZN(n646) );
  AND2_X1 U716 ( .A1(n646), .A2(n524), .ZN(n650) );
  NOR2_X1 U717 ( .A1(G299), .A2(n647), .ZN(n648) );
  XOR2_X1 U718 ( .A(KEYINPUT93), .B(n648), .Z(n649) );
  NOR2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT94), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n654), .B(KEYINPUT29), .ZN(n683) );
  XOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .Z(n937) );
  NOR2_X1 U723 ( .A1(n937), .A2(n655), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n656), .A2(G1961), .ZN(n657) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n661) );
  OR2_X1 U726 ( .A1(G301), .A2(n661), .ZN(n689) );
  AND2_X1 U727 ( .A1(G286), .A2(G8), .ZN(n660) );
  AND2_X1 U728 ( .A1(n689), .A2(n660), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n683), .A2(n659), .ZN(n680) );
  INV_X1 U730 ( .A(n660), .ZN(n670) );
  NAND2_X1 U731 ( .A1(n661), .A2(G301), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT95), .ZN(n668) );
  NOR2_X1 U733 ( .A1(G2084), .A2(n671), .ZN(n684) );
  NOR2_X1 U734 ( .A1(G1966), .A2(n713), .ZN(n663) );
  XNOR2_X1 U735 ( .A(KEYINPUT90), .B(n663), .ZN(n686) );
  NOR2_X1 U736 ( .A1(n684), .A2(n686), .ZN(n664) );
  NAND2_X1 U737 ( .A1(G8), .A2(n664), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT30), .B(n665), .ZN(n666) );
  NOR2_X1 U739 ( .A1(n666), .A2(G168), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT31), .B(n669), .Z(n691) );
  INV_X1 U742 ( .A(G8), .ZN(n676) );
  NOR2_X1 U743 ( .A1(G1971), .A2(n713), .ZN(n673) );
  NOR2_X1 U744 ( .A1(G2090), .A2(n671), .ZN(n672) );
  NOR2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n674), .A2(G303), .ZN(n675) );
  OR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(n681), .ZN(n696) );
  NAND2_X1 U750 ( .A1(G8), .A2(n684), .ZN(n685) );
  XNOR2_X1 U751 ( .A(KEYINPUT89), .B(n685), .ZN(n687) );
  OR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n692) );
  INV_X1 U753 ( .A(n692), .ZN(n688) );
  AND2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U755 ( .A1(n683), .A2(n690), .ZN(n694) );
  OR2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  AND2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n710) );
  NOR2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n964) );
  NOR2_X1 U760 ( .A1(G1971), .A2(G303), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n964), .A2(n697), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n710), .A2(n698), .ZN(n701) );
  NAND2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NAND2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n703) );
  INV_X1 U765 ( .A(KEYINPUT33), .ZN(n702) );
  NAND2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n964), .A2(KEYINPUT33), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n704), .A2(n713), .ZN(n706) );
  XOR2_X1 U769 ( .A(G1981), .B(G305), .Z(n953) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n709), .B(KEYINPUT96), .ZN(n716) );
  NOR2_X1 U773 ( .A1(G2090), .A2(G303), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G8), .A2(n711), .ZN(n712) );
  NAND2_X1 U775 ( .A1(n710), .A2(n712), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U778 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n719), .A2(n720), .ZN(n754) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n771) );
  NAND2_X1 U781 ( .A1(G104), .A2(n723), .ZN(n726) );
  BUF_X1 U782 ( .A(n724), .Z(n874) );
  NAND2_X1 U783 ( .A1(G140), .A2(n874), .ZN(n725) );
  NAND2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U785 ( .A(KEYINPUT34), .B(n727), .ZN(n732) );
  NAND2_X1 U786 ( .A1(G128), .A2(n888), .ZN(n729) );
  NAND2_X1 U787 ( .A1(G116), .A2(n889), .ZN(n728) );
  NAND2_X1 U788 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U789 ( .A(n730), .B(KEYINPUT35), .Z(n731) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U791 ( .A(KEYINPUT36), .B(n733), .Z(n734) );
  XNOR2_X1 U792 ( .A(KEYINPUT85), .B(n734), .ZN(n905) );
  XNOR2_X1 U793 ( .A(G2067), .B(KEYINPUT37), .ZN(n768) );
  NOR2_X1 U794 ( .A1(n905), .A2(n768), .ZN(n1021) );
  NAND2_X1 U795 ( .A1(n771), .A2(n1021), .ZN(n766) );
  NAND2_X1 U796 ( .A1(G105), .A2(n723), .ZN(n735) );
  XNOR2_X1 U797 ( .A(n735), .B(KEYINPUT38), .ZN(n742) );
  NAND2_X1 U798 ( .A1(G141), .A2(n874), .ZN(n737) );
  NAND2_X1 U799 ( .A1(G129), .A2(n888), .ZN(n736) );
  NAND2_X1 U800 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U801 ( .A1(G117), .A2(n889), .ZN(n738) );
  XNOR2_X1 U802 ( .A(KEYINPUT87), .B(n738), .ZN(n739) );
  NOR2_X1 U803 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U804 ( .A1(n742), .A2(n741), .ZN(n882) );
  NAND2_X1 U805 ( .A1(G1996), .A2(n882), .ZN(n751) );
  NAND2_X1 U806 ( .A1(G119), .A2(n888), .ZN(n744) );
  NAND2_X1 U807 ( .A1(G107), .A2(n889), .ZN(n743) );
  NAND2_X1 U808 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U809 ( .A1(n723), .A2(G95), .ZN(n745) );
  XOR2_X1 U810 ( .A(KEYINPUT86), .B(n745), .Z(n746) );
  NOR2_X1 U811 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U812 ( .A1(n874), .A2(G131), .ZN(n748) );
  NAND2_X1 U813 ( .A1(n749), .A2(n748), .ZN(n883) );
  NAND2_X1 U814 ( .A1(G1991), .A2(n883), .ZN(n750) );
  NAND2_X1 U815 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U816 ( .A(KEYINPUT88), .B(n752), .ZN(n1011) );
  NAND2_X1 U817 ( .A1(n771), .A2(n1011), .ZN(n761) );
  NAND2_X1 U818 ( .A1(n766), .A2(n761), .ZN(n753) );
  NOR2_X1 U819 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U820 ( .A(n755), .B(KEYINPUT98), .ZN(n757) );
  XNOR2_X1 U821 ( .A(G1986), .B(G290), .ZN(n961) );
  NAND2_X1 U822 ( .A1(n961), .A2(n771), .ZN(n756) );
  NAND2_X1 U823 ( .A1(n757), .A2(n756), .ZN(n774) );
  NOR2_X1 U824 ( .A1(G1996), .A2(n882), .ZN(n1007) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n759) );
  NOR2_X1 U826 ( .A1(G1991), .A2(n883), .ZN(n758) );
  XOR2_X1 U827 ( .A(KEYINPUT99), .B(n758), .Z(n1018) );
  NOR2_X1 U828 ( .A1(n759), .A2(n1018), .ZN(n760) );
  XOR2_X1 U829 ( .A(KEYINPUT100), .B(n760), .Z(n762) );
  NAND2_X1 U830 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U831 ( .A(KEYINPUT101), .B(n763), .ZN(n764) );
  NOR2_X1 U832 ( .A1(n1007), .A2(n764), .ZN(n765) );
  XNOR2_X1 U833 ( .A(KEYINPUT39), .B(n765), .ZN(n767) );
  NAND2_X1 U834 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U835 ( .A1(n905), .A2(n768), .ZN(n769) );
  XNOR2_X1 U836 ( .A(KEYINPUT102), .B(n769), .ZN(n1023) );
  NAND2_X1 U837 ( .A1(n770), .A2(n1023), .ZN(n772) );
  NAND2_X1 U838 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U839 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U840 ( .A(n775), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U842 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n777) );
  NAND2_X1 U843 ( .A1(G123), .A2(n888), .ZN(n776) );
  XNOR2_X1 U844 ( .A(n777), .B(n776), .ZN(n784) );
  NAND2_X1 U845 ( .A1(G99), .A2(n723), .ZN(n779) );
  NAND2_X1 U846 ( .A1(G135), .A2(n874), .ZN(n778) );
  NAND2_X1 U847 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U848 ( .A1(n889), .A2(G111), .ZN(n780) );
  XOR2_X1 U849 ( .A(KEYINPUT78), .B(n780), .Z(n781) );
  NOR2_X1 U850 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U851 ( .A1(n784), .A2(n783), .ZN(n1015) );
  XNOR2_X1 U852 ( .A(G2096), .B(n1015), .ZN(n785) );
  OR2_X1 U853 ( .A1(G2100), .A2(n785), .ZN(G156) );
  INV_X1 U854 ( .A(G120), .ZN(G236) );
  INV_X1 U855 ( .A(G69), .ZN(G235) );
  INV_X1 U856 ( .A(G108), .ZN(G238) );
  NAND2_X1 U857 ( .A1(G7), .A2(G661), .ZN(n786) );
  XNOR2_X1 U858 ( .A(n786), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U859 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n788) );
  XNOR2_X1 U860 ( .A(G223), .B(KEYINPUT69), .ZN(n839) );
  NAND2_X1 U861 ( .A1(G567), .A2(n839), .ZN(n787) );
  XNOR2_X1 U862 ( .A(n788), .B(n787), .ZN(G234) );
  INV_X1 U863 ( .A(G860), .ZN(n810) );
  OR2_X1 U864 ( .A1(n789), .A2(n810), .ZN(G153) );
  NAND2_X1 U865 ( .A1(G868), .A2(G301), .ZN(n791) );
  OR2_X1 U866 ( .A1(n951), .A2(G868), .ZN(n790) );
  NAND2_X1 U867 ( .A1(n791), .A2(n790), .ZN(G284) );
  NAND2_X1 U868 ( .A1(G868), .A2(G286), .ZN(n793) );
  INV_X1 U869 ( .A(G868), .ZN(n821) );
  NAND2_X1 U870 ( .A1(G299), .A2(n821), .ZN(n792) );
  NAND2_X1 U871 ( .A1(n793), .A2(n792), .ZN(G297) );
  NAND2_X1 U872 ( .A1(n810), .A2(G559), .ZN(n794) );
  NAND2_X1 U873 ( .A1(n794), .A2(n951), .ZN(n795) );
  XNOR2_X1 U874 ( .A(n795), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U875 ( .A1(G868), .A2(n789), .ZN(n798) );
  NAND2_X1 U876 ( .A1(G868), .A2(n951), .ZN(n796) );
  NOR2_X1 U877 ( .A1(G559), .A2(n796), .ZN(n797) );
  NOR2_X1 U878 ( .A1(n798), .A2(n797), .ZN(G282) );
  NAND2_X1 U879 ( .A1(G93), .A2(n523), .ZN(n802) );
  NAND2_X1 U880 ( .A1(G67), .A2(n800), .ZN(n801) );
  NAND2_X1 U881 ( .A1(n802), .A2(n801), .ZN(n808) );
  NAND2_X1 U882 ( .A1(G80), .A2(n803), .ZN(n806) );
  NAND2_X1 U883 ( .A1(G55), .A2(n804), .ZN(n805) );
  NAND2_X1 U884 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U885 ( .A1(n808), .A2(n807), .ZN(n822) );
  NAND2_X1 U886 ( .A1(G559), .A2(n951), .ZN(n809) );
  XOR2_X1 U887 ( .A(n789), .B(n809), .Z(n819) );
  NAND2_X1 U888 ( .A1(n810), .A2(n819), .ZN(n811) );
  XNOR2_X1 U889 ( .A(n811), .B(KEYINPUT79), .ZN(n812) );
  XOR2_X1 U890 ( .A(n822), .B(n812), .Z(G145) );
  INV_X1 U891 ( .A(G303), .ZN(G166) );
  XOR2_X1 U892 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n813) );
  XNOR2_X1 U893 ( .A(G288), .B(n813), .ZN(n816) );
  XNOR2_X1 U894 ( .A(G166), .B(G290), .ZN(n814) );
  XNOR2_X1 U895 ( .A(n814), .B(G299), .ZN(n815) );
  XNOR2_X1 U896 ( .A(n816), .B(n815), .ZN(n818) );
  XOR2_X1 U897 ( .A(G305), .B(n822), .Z(n817) );
  XNOR2_X1 U898 ( .A(n818), .B(n817), .ZN(n908) );
  XOR2_X1 U899 ( .A(n908), .B(n819), .Z(n820) );
  NOR2_X1 U900 ( .A1(n821), .A2(n820), .ZN(n824) );
  NOR2_X1 U901 ( .A1(G868), .A2(n822), .ZN(n823) );
  NOR2_X1 U902 ( .A1(n824), .A2(n823), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2078), .A2(G2084), .ZN(n825) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n825), .Z(n826) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n826), .ZN(n827) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n827), .ZN(n828) );
  NAND2_X1 U907 ( .A1(n828), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U909 ( .A1(G235), .A2(G236), .ZN(n829) );
  XOR2_X1 U910 ( .A(KEYINPUT84), .B(n829), .Z(n830) );
  NOR2_X1 U911 ( .A1(G238), .A2(n830), .ZN(n831) );
  NAND2_X1 U912 ( .A1(G57), .A2(n831), .ZN(n845) );
  NAND2_X1 U913 ( .A1(n845), .A2(G567), .ZN(n837) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n833) );
  NAND2_X1 U915 ( .A1(G132), .A2(G82), .ZN(n832) );
  XNOR2_X1 U916 ( .A(n833), .B(n832), .ZN(n834) );
  NOR2_X1 U917 ( .A1(n834), .A2(G218), .ZN(n835) );
  NAND2_X1 U918 ( .A1(G96), .A2(n835), .ZN(n846) );
  NAND2_X1 U919 ( .A1(n846), .A2(G2106), .ZN(n836) );
  NAND2_X1 U920 ( .A1(n837), .A2(n836), .ZN(n847) );
  NAND2_X1 U921 ( .A1(G483), .A2(G661), .ZN(n838) );
  NOR2_X1 U922 ( .A1(n847), .A2(n838), .ZN(n844) );
  NAND2_X1 U923 ( .A1(n844), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n839), .ZN(G217) );
  INV_X1 U925 ( .A(G661), .ZN(n841) );
  NAND2_X1 U926 ( .A1(G2), .A2(G15), .ZN(n840) );
  NOR2_X1 U927 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U928 ( .A(KEYINPUT106), .B(n842), .Z(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U930 ( .A1(n844), .A2(n843), .ZN(G188) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  NOR2_X1 U935 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n847), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2084), .Z(n849) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2078), .ZN(n848) );
  XNOR2_X1 U940 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U941 ( .A(n850), .B(G2100), .Z(n852) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2090), .ZN(n851) );
  XNOR2_X1 U943 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U944 ( .A(G2096), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U945 ( .A(G2678), .B(KEYINPUT107), .ZN(n853) );
  XNOR2_X1 U946 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U947 ( .A(n856), .B(n855), .Z(G227) );
  XNOR2_X1 U948 ( .A(G1991), .B(KEYINPUT108), .ZN(n866) );
  XOR2_X1 U949 ( .A(G1976), .B(G1961), .Z(n858) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1986), .ZN(n857) );
  XNOR2_X1 U951 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U952 ( .A(G1971), .B(G1956), .Z(n860) );
  XNOR2_X1 U953 ( .A(G1981), .B(G1966), .ZN(n859) );
  XNOR2_X1 U954 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U955 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT41), .ZN(n863) );
  XNOR2_X1 U957 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U958 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n888), .ZN(n867) );
  XNOR2_X1 U960 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U961 ( .A1(n723), .A2(G100), .ZN(n868) );
  NAND2_X1 U962 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U963 ( .A1(G136), .A2(n874), .ZN(n871) );
  NAND2_X1 U964 ( .A1(G112), .A2(n889), .ZN(n870) );
  NAND2_X1 U965 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U966 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G103), .A2(n723), .ZN(n876) );
  NAND2_X1 U968 ( .A1(G139), .A2(n874), .ZN(n875) );
  NAND2_X1 U969 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U970 ( .A1(G127), .A2(n888), .ZN(n878) );
  NAND2_X1 U971 ( .A1(G115), .A2(n889), .ZN(n877) );
  NAND2_X1 U972 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U974 ( .A1(n881), .A2(n880), .ZN(n1000) );
  XNOR2_X1 U975 ( .A(n1000), .B(n882), .ZN(n884) );
  XNOR2_X1 U976 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U977 ( .A(G160), .B(n885), .ZN(n904) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n887) );
  XNOR2_X1 U979 ( .A(n1015), .B(KEYINPUT111), .ZN(n886) );
  XNOR2_X1 U980 ( .A(n887), .B(n886), .ZN(n900) );
  NAND2_X1 U981 ( .A1(G130), .A2(n888), .ZN(n891) );
  NAND2_X1 U982 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U983 ( .A1(n891), .A2(n890), .ZN(n898) );
  XNOR2_X1 U984 ( .A(KEYINPUT110), .B(KEYINPUT45), .ZN(n896) );
  NAND2_X1 U985 ( .A1(n874), .A2(G142), .ZN(n894) );
  NAND2_X1 U986 ( .A1(n723), .A2(G106), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT109), .B(n892), .Z(n893) );
  NAND2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U990 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U991 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U992 ( .A(G164), .B(G162), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U994 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U995 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U996 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U997 ( .A(n908), .B(n789), .ZN(n909) );
  XNOR2_X1 U998 ( .A(n909), .B(G286), .ZN(n911) );
  XOR2_X1 U999 ( .A(n951), .B(G171), .Z(n910) );
  XNOR2_X1 U1000 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n912), .ZN(G397) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2443), .Z(n914) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2446), .ZN(n913) );
  XNOR2_X1 U1004 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1005 ( .A(n915), .B(G2430), .Z(n917) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n916) );
  XNOR2_X1 U1007 ( .A(n917), .B(n916), .ZN(n921) );
  XOR2_X1 U1008 ( .A(KEYINPUT105), .B(G2435), .Z(n919) );
  XNOR2_X1 U1009 ( .A(KEYINPUT104), .B(G2438), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1011 ( .A(n921), .B(n920), .Z(n923) );
  XNOR2_X1 U1012 ( .A(G2427), .B(KEYINPUT103), .ZN(n922) );
  XNOR2_X1 U1013 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1014 ( .A1(n924), .A2(G14), .ZN(n930) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1020 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G57), .ZN(G237) );
  INV_X1 U1023 ( .A(n930), .ZN(G401) );
  XNOR2_X1 U1024 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1039) );
  XOR2_X1 U1025 ( .A(G1991), .B(G25), .Z(n931) );
  NAND2_X1 U1026 ( .A1(n931), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1027 ( .A(G2067), .B(G26), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(G33), .B(G2072), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(n934), .B(KEYINPUT119), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(G1996), .B(G32), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G27), .B(n937), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT53), .B(n942), .ZN(n946) );
  XOR2_X1 U1037 ( .A(KEYINPUT120), .B(G34), .Z(n944) );
  XNOR2_X1 U1038 ( .A(G2084), .B(KEYINPUT54), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n944), .B(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G35), .B(G2090), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1043 ( .A(KEYINPUT55), .B(n949), .Z(n950) );
  NOR2_X1 U1044 ( .A1(G29), .A2(n950), .ZN(n1037) );
  XOR2_X1 U1045 ( .A(KEYINPUT56), .B(G16), .Z(n975) );
  XNOR2_X1 U1046 ( .A(n951), .B(G1348), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n952), .B(KEYINPUT121), .ZN(n973) );
  XNOR2_X1 U1048 ( .A(G171), .B(G1961), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G168), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n955), .B(KEYINPUT57), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G1341), .B(n789), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n971) );
  XNOR2_X1 U1055 ( .A(G166), .B(G1971), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G1956), .B(G299), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n969) );
  INV_X1 U1059 ( .A(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT122), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n1034) );
  XNOR2_X1 U1066 ( .A(G1348), .B(KEYINPUT59), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n976), .B(G4), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G19), .B(G1341), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G20), .B(G1956), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1074 ( .A(KEYINPUT60), .B(n983), .Z(n985) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n986), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G1961), .B(KEYINPUT123), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(G5), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n996) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(G23), .B(G1976), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1084 ( .A(G1986), .B(G24), .Z(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT58), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT61), .B(n997), .Z(n998) );
  NOR2_X1 U1089 ( .A1(G16), .A2(n998), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT125), .B(n999), .ZN(n1032) );
  XOR2_X1 U1091 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n1005) );
  XOR2_X1 U1092 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(n1003), .B(KEYINPUT50), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(n1005), .B(n1004), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT115), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(KEYINPUT51), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1026) );
  XNOR2_X1 U1103 ( .A(G160), .B(G2084), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(n1014), .B(KEYINPUT112), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1019), .B(KEYINPUT113), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT114), .B(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1027), .Z(n1028) );
  NOR2_X1 U1113 ( .A1(KEYINPUT55), .A2(n1028), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(KEYINPUT118), .B(n1029), .Z(n1030) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1035), .A2(G11), .ZN(n1036) );
  NOR2_X1 U1119 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1120 ( .A(n1039), .B(n1038), .ZN(G311) );
  XNOR2_X1 U1121 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

