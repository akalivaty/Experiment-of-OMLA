

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U326 ( .A(KEYINPUT96), .B(n466), .ZN(n536) );
  NOR2_X1 U327 ( .A1(n468), .A2(n517), .ZN(n469) );
  XNOR2_X1 U328 ( .A(n354), .B(n353), .ZN(n554) );
  XNOR2_X2 U329 ( .A(KEYINPUT107), .B(n491), .ZN(n496) );
  NOR2_X1 U330 ( .A1(n536), .A2(n453), .ZN(n551) );
  XOR2_X1 U331 ( .A(n415), .B(n414), .Z(n294) );
  XNOR2_X1 U332 ( .A(n416), .B(n294), .ZN(n417) );
  XNOR2_X1 U333 ( .A(n418), .B(n417), .ZN(n422) );
  INV_X1 U334 ( .A(G218GAT), .ZN(n456) );
  NOR2_X1 U335 ( .A1(n460), .A2(n454), .ZN(n585) );
  XOR2_X1 U336 ( .A(n428), .B(KEYINPUT41), .Z(n561) );
  XNOR2_X1 U337 ( .A(n456), .B(KEYINPUT62), .ZN(n457) );
  XNOR2_X1 U338 ( .A(n458), .B(n457), .ZN(G1355GAT) );
  XNOR2_X1 U339 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n295), .B(G29GAT), .ZN(n296) );
  XOR2_X1 U341 ( .A(n296), .B(KEYINPUT8), .Z(n298) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G50GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n393) );
  XOR2_X1 U344 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n300) );
  XNOR2_X1 U345 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n393), .B(n301), .ZN(n311) );
  XOR2_X1 U348 ( .A(KEYINPUT65), .B(KEYINPUT79), .Z(n303) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .Z(n408) );
  XOR2_X1 U352 ( .A(n408), .B(G162GAT), .Z(n305) );
  XOR2_X1 U353 ( .A(G190GAT), .B(G134GAT), .Z(n346) );
  XNOR2_X1 U354 ( .A(n346), .B(G218GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U356 ( .A(n307), .B(n306), .Z(n309) );
  NAND2_X1 U357 ( .A1(G232GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U359 ( .A(n311), .B(n310), .Z(n548) );
  XOR2_X1 U360 ( .A(KEYINPUT36), .B(n548), .Z(n485) );
  XOR2_X1 U361 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n313) );
  XNOR2_X1 U362 ( .A(G78GAT), .B(KEYINPUT93), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U364 ( .A(KEYINPUT91), .B(G162GAT), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(n316), .ZN(n372) );
  XNOR2_X1 U368 ( .A(n317), .B(n372), .ZN(n325) );
  XOR2_X1 U369 ( .A(G148GAT), .B(G155GAT), .Z(n319) );
  XNOR2_X1 U370 ( .A(G22GAT), .B(G211GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U372 ( .A(KEYINPUT24), .B(G204GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(KEYINPUT78), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n327) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U380 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U381 ( .A(KEYINPUT21), .B(G218GAT), .Z(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(G197GAT), .B(n332), .Z(n439) );
  XOR2_X1 U385 ( .A(G106GAT), .B(KEYINPUT73), .Z(n415) );
  XNOR2_X1 U386 ( .A(n439), .B(n415), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n552) );
  XOR2_X1 U388 ( .A(G176GAT), .B(KEYINPUT85), .Z(n336) );
  XNOR2_X1 U389 ( .A(G127GAT), .B(G120GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n354) );
  XOR2_X1 U391 ( .A(G113GAT), .B(KEYINPUT0), .Z(n359) );
  XNOR2_X1 U392 ( .A(G43GAT), .B(n359), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n337), .B(G99GAT), .ZN(n341) );
  XOR2_X1 U394 ( .A(G183GAT), .B(G71GAT), .Z(n339) );
  XNOR2_X1 U395 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U397 ( .A(n341), .B(n340), .Z(n352) );
  XOR2_X1 U398 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n343) );
  XNOR2_X1 U399 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n350) );
  XOR2_X1 U401 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n345) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n440) );
  XOR2_X1 U404 ( .A(n346), .B(n440), .Z(n348) );
  NAND2_X1 U405 ( .A1(G227GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n353) );
  NOR2_X1 U409 ( .A1(n552), .A2(n554), .ZN(n356) );
  XNOR2_X1 U410 ( .A(KEYINPUT26), .B(KEYINPUT103), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n460) );
  XOR2_X1 U412 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n371) );
  XOR2_X1 U415 ( .A(G120GAT), .B(G148GAT), .Z(n409) );
  XOR2_X1 U416 ( .A(G85GAT), .B(n409), .Z(n361) );
  XNOR2_X1 U417 ( .A(G134GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U419 ( .A(n362), .B(KEYINPUT94), .Z(n369) );
  XOR2_X1 U420 ( .A(G57GAT), .B(G155GAT), .Z(n364) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(G127GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n387) );
  XOR2_X1 U423 ( .A(n387), .B(KEYINPUT95), .Z(n366) );
  NAND2_X1 U424 ( .A1(G225GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(G29GAT), .B(n367), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n466) );
  INV_X1 U430 ( .A(n548), .ZN(n573) );
  XOR2_X1 U431 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n375) );
  NAND2_X1 U432 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U434 ( .A(n376), .B(KEYINPUT80), .Z(n380) );
  XNOR2_X1 U435 ( .A(G22GAT), .B(G15GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n377), .B(KEYINPUT69), .ZN(n394) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(G183GAT), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n378), .B(G211GAT), .ZN(n438) );
  XNOR2_X1 U439 ( .A(n394), .B(n438), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n382) );
  XNOR2_X1 U442 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U444 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U445 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n386) );
  XNOR2_X1 U446 ( .A(G71GAT), .B(G78GAT), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n405) );
  XNOR2_X1 U448 ( .A(n387), .B(n405), .ZN(n388) );
  XOR2_X1 U449 ( .A(n389), .B(n388), .Z(n584) );
  XNOR2_X1 U450 ( .A(n584), .B(KEYINPUT112), .ZN(n566) );
  XOR2_X1 U451 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n391) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n404) );
  XOR2_X1 U455 ( .A(G197GAT), .B(G141GAT), .Z(n396) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(n394), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U458 ( .A(G8GAT), .B(KEYINPUT68), .Z(n398) );
  NAND2_X1 U459 ( .A1(G229GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U461 ( .A(n400), .B(n399), .Z(n402) );
  XNOR2_X1 U462 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U464 ( .A(n404), .B(n403), .Z(n501) );
  XOR2_X1 U465 ( .A(n405), .B(KEYINPUT74), .Z(n407) );
  NAND2_X1 U466 ( .A1(G230GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n418) );
  XOR2_X1 U468 ( .A(KEYINPUT33), .B(n408), .Z(n411) );
  XNOR2_X1 U469 ( .A(G57GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n416) );
  XOR2_X1 U471 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U474 ( .A(G92GAT), .B(G64GAT), .Z(n420) );
  XNOR2_X1 U475 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U477 ( .A(G176GAT), .B(n421), .Z(n437) );
  XOR2_X1 U478 ( .A(n422), .B(n437), .Z(n581) );
  INV_X1 U479 ( .A(n581), .ZN(n428) );
  NOR2_X1 U480 ( .A1(n501), .A2(n561), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n423), .B(KEYINPUT46), .ZN(n424) );
  NOR2_X1 U482 ( .A1(n566), .A2(n424), .ZN(n425) );
  NAND2_X1 U483 ( .A1(n573), .A2(n425), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n426), .B(KEYINPUT47), .ZN(n433) );
  INV_X1 U485 ( .A(n584), .ZN(n487) );
  NOR2_X1 U486 ( .A1(n487), .A2(n485), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n427), .B(KEYINPUT45), .ZN(n429) );
  NAND2_X1 U488 ( .A1(n429), .A2(n428), .ZN(n431) );
  XOR2_X1 U489 ( .A(n501), .B(KEYINPUT71), .Z(n556) );
  INV_X1 U490 ( .A(n556), .ZN(n430) );
  NOR2_X1 U491 ( .A1(n431), .A2(n430), .ZN(n432) );
  NOR2_X1 U492 ( .A1(n433), .A2(n432), .ZN(n436) );
  XOR2_X1 U493 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n434) );
  XNOR2_X1 U494 ( .A(KEYINPUT48), .B(n434), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n538) );
  XOR2_X1 U496 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n450) );
  NAND2_X1 U499 ( .A1(G226GAT), .A2(G233GAT), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT97), .B(KEYINPUT100), .Z(n444) );
  XNOR2_X1 U501 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U503 ( .A(G36GAT), .B(G190GAT), .Z(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n514) );
  INV_X1 U507 ( .A(n514), .ZN(n451) );
  NOR2_X1 U508 ( .A1(n538), .A2(n451), .ZN(n452) );
  XOR2_X1 U509 ( .A(KEYINPUT54), .B(n452), .Z(n453) );
  INV_X1 U510 ( .A(n551), .ZN(n454) );
  INV_X1 U511 ( .A(n585), .ZN(n455) );
  NOR2_X1 U512 ( .A1(n485), .A2(n455), .ZN(n458) );
  NOR2_X1 U513 ( .A1(n581), .A2(n556), .ZN(n489) );
  XOR2_X1 U514 ( .A(KEYINPUT27), .B(KEYINPUT101), .Z(n459) );
  XOR2_X1 U515 ( .A(n514), .B(n459), .Z(n468) );
  NOR2_X1 U516 ( .A1(n460), .A2(n468), .ZN(n535) );
  NAND2_X1 U517 ( .A1(n514), .A2(n554), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n552), .A2(n461), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n535), .A2(n463), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT104), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n472) );
  XOR2_X1 U523 ( .A(n552), .B(KEYINPUT66), .Z(n467) );
  XNOR2_X1 U524 ( .A(KEYINPUT28), .B(n467), .ZN(n517) );
  NAND2_X1 U525 ( .A1(n536), .A2(n469), .ZN(n522) );
  NOR2_X1 U526 ( .A1(n554), .A2(n522), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT102), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT105), .B(n473), .Z(n484) );
  NAND2_X1 U530 ( .A1(n573), .A2(n584), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT16), .B(n474), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n484), .A2(n475), .ZN(n502) );
  AND2_X1 U533 ( .A1(n489), .A2(n502), .ZN(n482) );
  NAND2_X1 U534 ( .A1(n536), .A2(n482), .ZN(n476) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n482), .A2(n514), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n480) );
  NAND2_X1 U540 ( .A1(n482), .A2(n554), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n517), .A2(n482), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT39), .B(KEYINPUT108), .Z(n493) );
  NOR2_X1 U546 ( .A1(n485), .A2(n484), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n488), .ZN(n512) );
  NAND2_X1 U549 ( .A1(n489), .A2(n512), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT38), .ZN(n491) );
  NAND2_X1 U551 ( .A1(n536), .A2(n496), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n496), .A2(n514), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n554), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  XOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT109), .Z(n500) );
  NAND2_X1 U560 ( .A1(n496), .A2(n517), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  INV_X1 U562 ( .A(n501), .ZN(n576) );
  NOR2_X1 U563 ( .A1(n576), .A2(n561), .ZN(n511) );
  AND2_X1 U564 ( .A1(n511), .A2(n502), .ZN(n508) );
  NAND2_X1 U565 ( .A1(n508), .A2(n536), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(KEYINPUT110), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n514), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n554), .A2(n508), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n517), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  AND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n518) );
  NAND2_X1 U577 ( .A1(n536), .A2(n518), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n518), .A2(n514), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n554), .A2(n518), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n538), .A2(n522), .ZN(n523) );
  NAND2_X1 U588 ( .A1(n523), .A2(n554), .ZN(n531) );
  NOR2_X1 U589 ( .A1(n556), .A2(n531), .ZN(n524) );
  XOR2_X1 U590 ( .A(G113GAT), .B(n524), .Z(G1340GAT) );
  NOR2_X1 U591 ( .A1(n561), .A2(n531), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n529) );
  INV_X1 U595 ( .A(n531), .ZN(n527) );
  NAND2_X1 U596 ( .A1(n527), .A2(n566), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U598 ( .A(G127GAT), .B(n530), .Z(G1342GAT) );
  NOR2_X1 U599 ( .A1(n573), .A2(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U602 ( .A(G134GAT), .B(n534), .Z(G1343GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U604 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n549), .A2(n576), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XNOR2_X1 U609 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n546) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .Z(n544) );
  INV_X1 U611 ( .A(n561), .ZN(n542) );
  NAND2_X1 U612 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n584), .A2(n549), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT55), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n572) );
  NOR2_X1 U622 ( .A1(n556), .A2(n572), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT119), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n561), .A2(n572), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .Z(n569) );
  INV_X1 U633 ( .A(n572), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n575) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(n575), .B(n574), .Z(G1351GAT) );
  NAND2_X1 U641 ( .A1(n585), .A2(n576), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
endmodule

