//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G137), .A3(new_n461), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n470), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  AOI211_X1 g047(.A(new_n472), .B(new_n461), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n463), .B(new_n465), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(new_n461), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n467), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n461), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n478), .B(new_n482), .C1(new_n486), .C2(G124), .ZN(G162));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n466), .B2(new_n467), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n467), .C2(new_n466), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n503), .ZN(new_n511));
  AOI21_X1  g086(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(G88), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G50), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G166));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n509), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n501), .B1(new_n517), .B2(KEYINPUT71), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n508), .A2(new_n519), .A3(new_n509), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n510), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n522), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT72), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT72), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G651), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(G52), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n521), .A2(new_n535), .B1(G90), .B2(new_n524), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n499), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(G81), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n540), .B1(new_n524), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n521), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n518), .A2(new_n520), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n518), .A2(new_n554), .A3(G53), .A4(new_n520), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n523), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n524), .B2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n524), .A2(G87), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n518), .A2(G49), .A3(new_n520), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n511), .A2(G74), .A3(new_n512), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n524), .A2(G87), .B1(new_n566), .B2(G651), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n565), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G288));
  AND2_X1   g149(.A1(new_n504), .A2(G86), .ZN(new_n575));
  AND2_X1   g150(.A1(G48), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n517), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n523), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n524), .A2(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT76), .B(G47), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n499), .B2(new_n584), .C1(new_n551), .C2(new_n585), .ZN(G290));
  AOI22_X1  g161(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n499), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G54), .B2(new_n521), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n504), .A2(G92), .A3(new_n517), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G171), .B2(new_n593), .ZN(G284));
  OAI21_X1  g170(.A(new_n594), .B1(G171), .B2(new_n593), .ZN(G321));
  NOR2_X1   g171(.A1(G168), .A2(new_n593), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT77), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(G868), .B2(new_n599), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(G868), .B2(new_n599), .ZN(G280));
  INV_X1    g176(.A(new_n592), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n544), .A2(new_n593), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n592), .A2(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n593), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n464), .A2(new_n462), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n461), .A2(G111), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT78), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n613), .B2(KEYINPUT78), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n480), .A2(G135), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT69), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n485), .B(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G123), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n612), .A2(G2100), .B1(G2096), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n622), .B(new_n623), .C1(G2100), .C2(new_n612), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G1341), .ZN(new_n633));
  INV_X1    g208(.A(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n635), .A2(new_n639), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  INV_X1    g224(.A(new_n646), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n650), .B2(new_n644), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n644), .B(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n651), .B1(new_n653), .B2(new_n650), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n650), .A3(new_n647), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT82), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  MUX2_X1   g245(.A(new_n670), .B(new_n669), .S(new_n662), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(KEYINPUT94), .ZN(new_n679));
  MUX2_X1   g254(.A(G23), .B(new_n568), .S(G16), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G1971), .ZN(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(G1971), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n683), .A2(new_n688), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT34), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT34), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n480), .A2(G131), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n461), .A2(G107), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  INV_X1    g273(.A(G119), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n696), .B1(new_n697), .B2(new_n698), .C1(new_n619), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT84), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT83), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT83), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n701), .S(new_n705), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT85), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(G16), .A2(G24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G290), .B2(new_n684), .ZN(new_n711));
  INV_X1    g286(.A(G1986), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n713), .B(new_n714), .C1(KEYINPUT88), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n694), .A2(new_n695), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(KEYINPUT88), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT89), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n694), .A2(new_n695), .A3(new_n717), .A4(new_n720), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n705), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n705), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2090), .ZN(new_n728));
  NOR2_X1   g303(.A1(G5), .A2(G16), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G171), .B2(G16), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT93), .B(G1961), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n684), .A2(G4), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n602), .B2(new_n684), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(new_n634), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n684), .A2(G19), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT90), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n544), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1341), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n702), .A2(G32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n486), .A2(G129), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n462), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT26), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n744), .B(new_n746), .C1(new_n480), .C2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n702), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n684), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n684), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n751), .A2(new_n752), .B1(G1966), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G1966), .B2(new_n754), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT31), .B(G11), .Z(new_n757));
  INV_X1    g332(.A(new_n705), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n621), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT92), .B(G28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n757), .B(new_n759), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G164), .A2(new_n758), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G27), .B2(new_n758), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n764), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n702), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G139), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n479), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n464), .A2(G127), .ZN(new_n777));
  NAND2_X1  g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n461), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n771), .B1(new_n780), .B2(new_n702), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n751), .B2(new_n752), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n741), .A2(new_n756), .A3(new_n770), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n758), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n486), .A2(G128), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G116), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n480), .B2(G140), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G29), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(KEYINPUT91), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(KEYINPUT91), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2067), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n684), .A2(G20), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT23), .Z(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G299), .B2(G16), .ZN(new_n800));
  INV_X1    g375(.A(G1956), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G34), .ZN(new_n804));
  AOI22_X1  g379(.A1(G160), .A2(G29), .B1(new_n758), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G2084), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n733), .A2(new_n784), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n679), .B1(new_n724), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g385(.A(KEYINPUT94), .B(new_n808), .C1(new_n722), .C2(new_n723), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(G311));
  NAND2_X1  g387(.A1(new_n724), .A2(new_n809), .ZN(G150));
  NAND2_X1  g388(.A1(new_n524), .A2(G93), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n814), .B1(new_n499), .B2(new_n815), .C1(new_n816), .C2(new_n551), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT95), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n544), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n544), .A2(new_n817), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n602), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  AOI21_X1  g400(.A(G860), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n818), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(G145));
  XNOR2_X1  g405(.A(G160), .B(new_n621), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(G162), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n480), .A2(G142), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n461), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G130), .B2(new_n486), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(new_n610), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n700), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n748), .B(new_n792), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n495), .A2(new_n497), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n489), .A2(new_n490), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT96), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT96), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n840), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n780), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  INV_X1    g424(.A(new_n497), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n496), .B1(new_n464), .B2(new_n493), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n849), .B1(new_n852), .B2(new_n491), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT96), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n840), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n780), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n839), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n838), .B(new_n700), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n780), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n846), .A2(new_n847), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n832), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT97), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(KEYINPUT99), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(new_n839), .C1(new_n848), .C2(new_n857), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n865), .A2(new_n832), .A3(new_n862), .A4(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(G37), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n864), .A2(new_n870), .A3(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(G395));
  AND2_X1   g451(.A1(new_n819), .A2(new_n820), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n606), .ZN(new_n878));
  XOR2_X1   g453(.A(G299), .B(new_n592), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n821), .B(new_n606), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n879), .B(KEYINPUT41), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(G290), .B(G305), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n568), .B(G166), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n881), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n881), .B2(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n818), .A2(new_n593), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  XNOR2_X1  g469(.A(G295), .B(new_n894), .ZN(G331));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  OAI21_X1  g471(.A(G168), .B1(G301), .B2(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(G301), .A2(KEYINPUT103), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n897), .B(new_n898), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n821), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n897), .B(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n877), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n883), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n902), .A3(new_n879), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n887), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n887), .B1(new_n904), .B2(new_n905), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n896), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n880), .A2(new_n900), .A3(new_n902), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n911), .ZN(new_n914));
  INV_X1    g489(.A(new_n887), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n869), .A3(new_n906), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n910), .B1(new_n917), .B2(new_n896), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT44), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n908), .B2(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n465), .A2(G40), .A3(new_n463), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n472), .B1(new_n927), .B2(new_n461), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n470), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n925), .B(new_n930), .C1(new_n855), .C2(G1384), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n931), .A2(G1996), .A3(new_n748), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT105), .ZN(new_n933));
  INV_X1    g508(.A(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n792), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n749), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n933), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n700), .B(new_n708), .Z(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(G290), .B(G1986), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT125), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT111), .B(G1981), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n577), .A2(new_n581), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1981), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n577), .B2(new_n581), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n945), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n951), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT49), .A3(new_n948), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n841), .B2(new_n842), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n930), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1976), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n570), .A2(new_n572), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n571), .A2(G1976), .A3(new_n565), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n957), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n962), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT52), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n958), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n841), .A2(new_n842), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n925), .A2(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n930), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n977), .A3(new_n806), .A4(new_n930), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n955), .B(G286), .C1(new_n973), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n853), .A2(new_n854), .A3(new_n969), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT106), .B1(new_n956), .B2(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n925), .C1(G164), .C2(G1384), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n930), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n974), .A2(new_n930), .A3(new_n977), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n955), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT108), .B(KEYINPUT55), .Z(new_n992));
  OAI211_X1 g567(.A(G8), .B(new_n992), .C1(new_n507), .C2(new_n515), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n513), .A2(new_n514), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n517), .ZN(new_n995));
  INV_X1    g570(.A(G62), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n502), .B2(new_n503), .ZN(new_n997));
  INV_X1    g572(.A(new_n506), .ZN(new_n998));
  OAI21_X1  g573(.A(G651), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n955), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n993), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n991), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT63), .B1(new_n980), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G288), .A2(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n949), .B1(new_n1006), .B2(new_n958), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n957), .B(KEYINPUT112), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT63), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n968), .A2(new_n975), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n956), .A2(new_n976), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1012), .A2(new_n989), .A3(new_n930), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n955), .B1(new_n987), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1010), .B(new_n979), .C1(new_n1015), .C2(new_n1003), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1003), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n993), .B(KEYINPUT109), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT110), .B1(new_n991), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n985), .A2(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  NOR4_X1   g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1020), .A4(new_n955), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1016), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1009), .B1(new_n1026), .B2(new_n966), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n982), .A2(new_n984), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n465), .A2(G40), .A3(new_n463), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n471), .B2(new_n473), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n845), .B2(new_n969), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT115), .Z(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT116), .B1(new_n985), .B2(new_n1034), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1012), .A2(new_n930), .A3(new_n1013), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n801), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n556), .A2(new_n1041), .A3(new_n560), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n556), .B2(new_n560), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n556), .A2(KEYINPUT113), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1042), .A2(new_n1043), .B1(new_n1044), .B2(KEYINPUT57), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G299), .A2(KEYINPUT114), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n556), .B2(KEYINPUT113), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n556), .A2(new_n1041), .A3(new_n560), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1040), .B(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1011), .A2(new_n1030), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT117), .B1(new_n930), .B2(new_n956), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n935), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n974), .A2(new_n930), .A3(new_n977), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n634), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n592), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1055), .A2(KEYINPUT119), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n592), .A2(new_n1058), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1067), .A3(new_n1063), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1051), .A2(KEYINPUT61), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1052), .B1(new_n1011), .B2(new_n1030), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n930), .A2(KEYINPUT117), .A3(new_n956), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT58), .B(G1341), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT118), .B(G1996), .Z(new_n1074));
  OAI22_X1  g649(.A1(new_n1072), .A2(new_n1073), .B1(new_n985), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n545), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(KEYINPUT59), .A3(new_n545), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1040), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1050), .A2(new_n1037), .A3(new_n1039), .A4(new_n1036), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n592), .B2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1069), .A2(new_n1085), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n985), .B2(G2078), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n971), .A2(new_n972), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1056), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT121), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1099), .A3(G171), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1029), .B(KEYINPUT122), .C1(new_n461), .C2(new_n927), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n927), .A2(new_n461), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n926), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1102), .A2(new_n1092), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n855), .A2(G1384), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n981), .B(new_n1106), .C1(new_n1107), .C2(KEYINPUT45), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1090), .A2(new_n1108), .A3(new_n1095), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1101), .B1(new_n1109), .B2(G171), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1095), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1028), .A2(new_n1031), .A3(new_n767), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1089), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1113), .A2(KEYINPUT123), .A3(G301), .A4(new_n1108), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1098), .A2(new_n1100), .A3(new_n1110), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n1096), .B2(G171), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1113), .A2(KEYINPUT124), .A3(new_n1108), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  AOI21_X1  g695(.A(G301), .B1(new_n1109), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n973), .A2(G168), .A3(new_n978), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(G8), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G168), .B1(new_n973), .B2(new_n978), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(G8), .A3(new_n1125), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1128), .B1(new_n1131), .B2(KEYINPUT51), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n966), .B1(new_n1015), .B2(new_n1003), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1124), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1117), .A2(new_n1123), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n944), .B(new_n1027), .C1(new_n1088), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1125), .A2(G8), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT51), .B1(new_n1137), .B2(new_n1129), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1127), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1139), .B(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1022), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n991), .A2(KEYINPUT110), .A3(new_n1021), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1133), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1141), .A2(KEYINPUT126), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1142), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1132), .A2(new_n1140), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(KEYINPUT62), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1136), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1087), .A2(new_n1082), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1080), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1051), .B2(KEYINPUT61), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1081), .A2(new_n1082), .A3(KEYINPUT61), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1068), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1067), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1155), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  NOR4_X1   g737(.A1(new_n1122), .A2(new_n1124), .A3(new_n1133), .A4(new_n1132), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(new_n1117), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n944), .B1(new_n1164), .B2(new_n1027), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n943), .B1(new_n1154), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n931), .B1(new_n936), .B2(new_n749), .ZN(new_n1167));
  OR3_X1    g742(.A1(new_n931), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT46), .B1(new_n931), .B2(G1996), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1171));
  XNOR2_X1  g746(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n931), .A2(G1986), .A3(G290), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT48), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n941), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n701), .A2(new_n708), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n939), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n787), .A2(new_n935), .A3(new_n791), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n931), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1166), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g756(.A(G319), .ZN(new_n1183));
  OR2_X1    g757(.A1(G227), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G229), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1185), .B1(new_n642), .B2(new_n641), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1186), .B1(new_n864), .B2(new_n870), .ZN(new_n1187));
  AND2_X1   g761(.A1(new_n1187), .A2(new_n921), .ZN(G308));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n921), .ZN(G225));
endmodule


