//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n542, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132, new_n1133;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n472), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g054(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n475), .B1(new_n482), .B2(G2105), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n467), .A2(new_n470), .A3(G2105), .A4(new_n472), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n473), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(new_n470), .A3(new_n472), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n478), .B2(new_n479), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n504), .A2(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n505), .B2(KEYINPUT70), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(G88), .B1(new_n514), .B2(G50), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(G166));
  XOR2_X1   g091(.A(KEYINPUT71), .B(G89), .Z(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n512), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(G168));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(G77), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n502), .A2(new_n503), .ZN(new_n528));
  INV_X1    g103(.A(G64), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n526), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n532), .B1(new_n531), .B2(new_n530), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n513), .A2(G90), .B1(new_n514), .B2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  AOI22_X1  g111(.A1(new_n513), .A2(G81), .B1(new_n514), .B2(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(new_n513), .A2(G91), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n514), .A2(G53), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n549), .A2(KEYINPUT9), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(KEYINPUT9), .ZN(new_n551));
  OAI221_X1 g126(.A(new_n547), .B1(new_n526), .B2(new_n548), .C1(new_n550), .C2(new_n551), .ZN(G299));
  INV_X1    g127(.A(G168), .ZN(G286));
  INV_X1    g128(.A(G166), .ZN(G303));
  AND3_X1   g129(.A1(new_n504), .A2(new_n511), .A3(G87), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n504), .A2(G74), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n514), .B2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G288));
  NAND2_X1  g135(.A1(new_n504), .A2(G61), .ZN(new_n561));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n526), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n504), .A2(new_n511), .A3(G86), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n526), .ZN(new_n570));
  INV_X1    g145(.A(G85), .ZN(new_n571));
  INV_X1    g146(.A(G47), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n512), .A2(new_n571), .B1(new_n518), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  INV_X1    g150(.A(G868), .ZN(new_n576));
  NOR2_X1   g151(.A1(G301), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n504), .A2(new_n511), .A3(G92), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n528), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n577), .B1(new_n589), .B2(new_n576), .ZN(G284));
  AOI21_X1  g165(.A(new_n577), .B1(new_n589), .B2(new_n576), .ZN(G321));
  NAND2_X1  g166(.A1(G299), .A2(new_n576), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n576), .B2(G168), .ZN(G297));
  OAI21_X1  g168(.A(new_n592), .B1(new_n576), .B2(G168), .ZN(G280));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n589), .B1(new_n595), .B2(G860), .ZN(G148));
  OAI21_X1  g171(.A(KEYINPUT77), .B1(new_n540), .B2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n595), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  MUX2_X1   g174(.A(KEYINPUT77), .B(new_n597), .S(new_n599), .Z(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n489), .A2(G135), .ZN(new_n602));
  INV_X1    g177(.A(new_n486), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G123), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n471), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n602), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT81), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2096), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n469), .A2(G2104), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT68), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n465), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT80), .B(G2100), .Z(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n617), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n609), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2430), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n633), .ZN(G401));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT17), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2084), .B(G2090), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n639), .A2(new_n641), .ZN(new_n646));
  NOR3_X1   g221(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n645), .A2(new_n641), .A3(new_n639), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n640), .A2(new_n645), .A3(new_n642), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G22), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G166), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(G1971), .Z(new_n678));
  NOR2_X1   g253(.A1(G6), .A2(G16), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n567), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT32), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(G16), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT33), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n678), .A2(new_n683), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  INV_X1    g269(.A(G107), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G2105), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  INV_X1    g272(.A(G119), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n486), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n489), .A2(G131), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT89), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n675), .A2(G24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n574), .B2(new_n675), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n692), .A2(new_n693), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT36), .Z(new_n715));
  INV_X1    g290(.A(G21), .ZN(new_n716));
  AOI21_X1  g291(.A(KEYINPUT95), .B1(new_n675), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G168), .A2(G16), .ZN(new_n718));
  MUX2_X1   g293(.A(KEYINPUT95), .B(new_n717), .S(new_n718), .Z(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G1966), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT97), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(G1966), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT31), .B(G11), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT96), .B(G28), .Z(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT30), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n724), .B2(KEYINPUT30), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n675), .A2(G5), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G171), .B2(new_n675), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(G1961), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  INV_X1    g307(.A(new_n608), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n721), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT98), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  NOR2_X1   g312(.A1(G4), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n589), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1348), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n732), .A2(G35), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT99), .Z(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n732), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT29), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(G2090), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n732), .A2(G32), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT26), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(G105), .B2(new_n465), .ZN(new_n752));
  INV_X1    g327(.A(G129), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n486), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G141), .B2(new_n489), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n732), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT27), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1996), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n736), .A2(new_n737), .A3(new_n746), .A4(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  NAND2_X1  g335(.A1(G164), .A2(G29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G27), .B2(G29), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n730), .A2(G1961), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n675), .A2(G20), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT23), .Z(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT100), .B(G1956), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n489), .A2(G139), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n770));
  NAND3_X1  g345(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n614), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n769), .B(new_n772), .C1(new_n773), .C2(new_n471), .ZN(new_n774));
  MUX2_X1   g349(.A(G33), .B(new_n774), .S(G29), .Z(new_n775));
  OAI21_X1  g350(.A(new_n768), .B1(G2072), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n732), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  OR2_X1    g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n780));
  INV_X1    g355(.A(G128), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n486), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G140), .B2(new_n489), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(new_n732), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT93), .Z(new_n785));
  AOI211_X1 g360(.A(new_n763), .B(new_n776), .C1(G2067), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n675), .A2(G19), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT92), .Z(new_n788));
  INV_X1    g363(.A(new_n540), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1341), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G160), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2084), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n775), .A2(G2072), .B1(new_n760), .B2(new_n762), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n791), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n785), .ZN(new_n801));
  INV_X1    g376(.A(G2067), .ZN(new_n802));
  INV_X1    g377(.A(G2090), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n744), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n786), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n715), .A2(new_n759), .A3(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  AOI22_X1  g382(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n526), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n512), .A2(new_n810), .B1(new_n518), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n539), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n789), .B2(new_n813), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n589), .A2(G559), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n816), .B(new_n817), .Z(new_n818));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n819));
  AOI21_X1  g394(.A(G860), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n813), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(G145));
  XNOR2_X1  g399(.A(new_n704), .B(new_n617), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n603), .A2(G130), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n471), .A2(G118), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n489), .A2(new_n829), .A3(G142), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n489), .B2(G142), .ZN(new_n831));
  OAI221_X1 g406(.A(new_n826), .B1(new_n827), .B2(new_n828), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n825), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n500), .A2(new_n498), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n603), .A2(G126), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n492), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n783), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n774), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n755), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(new_n840), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(KEYINPUT103), .A3(new_n843), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n834), .A2(KEYINPUT103), .A3(new_n841), .ZN(new_n845));
  XNOR2_X1  g420(.A(G160), .B(KEYINPUT101), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G162), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n608), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n834), .B2(new_n841), .ZN(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n850), .B2(new_n843), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g428(.A(new_n598), .B(KEYINPUT104), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n815), .ZN(new_n855));
  XNOR2_X1  g430(.A(G299), .B(new_n585), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G288), .B(G290), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT106), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G166), .B(new_n567), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT42), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n861), .A2(new_n863), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n861), .B2(new_n863), .ZN(new_n874));
  OAI21_X1  g449(.A(G868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n813), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(G868), .B2(new_n876), .ZN(G295));
  OAI21_X1  g452(.A(new_n875), .B1(G868), .B2(new_n876), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n879));
  AOI21_X1  g454(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n880));
  NOR2_X1   g455(.A1(G301), .A2(KEYINPUT107), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(new_n815), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n856), .ZN(new_n884));
  INV_X1    g459(.A(new_n871), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n882), .B(new_n815), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n860), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n885), .B1(new_n884), .B2(new_n887), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n879), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n862), .A2(new_n857), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n862), .B2(new_n859), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n884), .B1(new_n883), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n871), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n889), .A3(new_n888), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n892), .B1(new_n897), .B2(new_n879), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT44), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n896), .A2(new_n879), .A3(new_n889), .A4(new_n888), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n890), .B2(new_n891), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(G397));
  INV_X1    g480(.A(new_n475), .ZN(new_n906));
  INV_X1    g481(.A(new_n481), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n614), .B2(G125), .ZN(new_n908));
  OAI211_X1 g483(.A(G40), .B(new_n906), .C1(new_n908), .C2(new_n471), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n482), .A2(G2105), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n912), .A2(KEYINPUT108), .A3(G40), .A4(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(G164), .B2(G1384), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n704), .A2(new_n707), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n704), .A2(new_n707), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n755), .B(G1996), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n783), .B(G2067), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n574), .B(G1986), .Z(new_n924));
  OAI21_X1  g499(.A(new_n917), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(G164), .B2(G1384), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n614), .A2(new_n499), .B1(KEYINPUT4), .B2(new_n497), .ZN(new_n929));
  OAI211_X1 g504(.A(KEYINPUT112), .B(new_n928), .C1(new_n929), .C2(new_n494), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT108), .B1(G160), .B2(G40), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n934));
  INV_X1    g509(.A(G40), .ZN(new_n935));
  NOR4_X1   g510(.A1(new_n934), .A2(new_n910), .A3(new_n935), .A4(new_n475), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n837), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n932), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT121), .B(G1961), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n927), .A2(new_n944), .A3(new_n930), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n911), .A2(new_n913), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT122), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n941), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n938), .A2(new_n916), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n937), .A2(new_n955), .A3(KEYINPUT109), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n911), .A2(new_n938), .A3(new_n913), .A4(new_n916), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G2078), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(KEYINPUT53), .ZN(new_n961));
  AOI21_X1  g536(.A(G301), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  INV_X1    g538(.A(G2084), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n937), .A2(new_n964), .A3(new_n945), .A4(new_n947), .ZN(new_n965));
  INV_X1    g540(.A(G1966), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n911), .A2(new_n913), .A3(new_n938), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(new_n931), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n963), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G286), .A2(G8), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT120), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n969), .A2(KEYINPUT51), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n968), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n973), .B2(G8), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n973), .B2(new_n971), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n962), .B1(new_n978), .B2(KEYINPUT62), .ZN(new_n979));
  NOR2_X1   g554(.A1(G166), .A2(new_n963), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT55), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT110), .B(G1971), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n956), .A2(new_n959), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n837), .A2(new_n944), .A3(new_n928), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n911), .A2(new_n913), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n944), .B1(new_n927), .B2(new_n930), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n985), .A2(new_n986), .A3(G2090), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n981), .B1(new_n988), .B2(G8), .ZN(new_n989));
  OAI21_X1  g564(.A(G1981), .B1(new_n563), .B2(new_n566), .ZN(new_n990));
  INV_X1    g565(.A(G61), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n502), .B2(new_n503), .ZN(new_n992));
  INV_X1    g567(.A(new_n562), .ZN(new_n993));
  OAI21_X1  g568(.A(G651), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(new_n682), .A3(new_n564), .A4(new_n565), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n990), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n996), .A2(new_n997), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n911), .A2(new_n913), .A3(new_n927), .A4(new_n930), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(G8), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n685), .A2(G1976), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .A4(G8), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1004), .A3(G8), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1009), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT113), .B1(new_n1009), .B2(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n989), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n983), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n937), .A2(new_n803), .A3(new_n945), .A4(new_n947), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n956), .A2(new_n959), .A3(KEYINPUT111), .A4(new_n982), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(G8), .A3(new_n981), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT124), .B1(new_n979), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT124), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n974), .A2(new_n976), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n973), .A2(new_n971), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT51), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n974), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1022), .A2(new_n1023), .A3(new_n962), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1021), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n589), .A2(KEYINPUT60), .ZN(new_n1033));
  INV_X1    g608(.A(G1348), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n946), .B2(new_n948), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n937), .A2(new_n802), .A3(new_n927), .A4(new_n930), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n589), .A2(KEYINPUT60), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(new_n1036), .A3(KEYINPUT60), .A4(new_n589), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT58), .B(G1341), .Z(new_n1043));
  AND2_X1   g618(.A1(new_n1002), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT117), .B(G1996), .Z(new_n1045));
  NOR2_X1   g620(.A1(new_n957), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n540), .B(new_n1042), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n957), .A2(new_n1045), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1002), .A2(new_n1043), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n789), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1047), .B(KEYINPUT119), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  INV_X1    g628(.A(G1956), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n985), .B2(new_n986), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(G299), .B(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n937), .A2(new_n955), .A3(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1055), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1060), .B2(new_n1055), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1053), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1050), .A2(new_n1064), .A3(new_n1042), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1041), .A2(new_n1052), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1061), .A2(new_n1053), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT116), .B1(new_n1068), .B2(new_n1058), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1037), .A2(new_n589), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1069), .A2(new_n1073), .A3(new_n1071), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1066), .A2(new_n1072), .B1(new_n1074), .B2(new_n1061), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n954), .A2(new_n961), .A3(G301), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n909), .A2(KEYINPUT123), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n939), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n955), .B(new_n1079), .C1(KEYINPUT123), .C2(new_n909), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1080), .A2(new_n949), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(KEYINPUT53), .B2(new_n960), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1077), .B1(new_n1082), .B2(G171), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1027), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1081), .B(G301), .C1(KEYINPUT53), .C2(new_n960), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1077), .B1(new_n962), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1075), .A2(new_n1084), .A3(new_n1022), .A4(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n969), .A2(G168), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1013), .A2(new_n1019), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(KEYINPUT63), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(new_n1012), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1018), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(new_n981), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1097), .A3(new_n1019), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1019), .A2(new_n1012), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1002), .A2(G8), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1003), .A2(new_n1005), .A3(new_n685), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n995), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1088), .A2(new_n1099), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n925), .B1(new_n1032), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n917), .ZN(new_n1107));
  OR3_X1    g682(.A1(new_n1107), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT46), .B1(new_n1107), .B2(G1996), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n921), .A2(new_n755), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1108), .A2(new_n1109), .B1(new_n917), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT47), .Z(new_n1112));
  AND2_X1   g687(.A1(new_n923), .A2(new_n917), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT127), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1107), .A2(G1986), .A3(G290), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT48), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1112), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n922), .A2(new_n917), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1121), .A2(new_n919), .B1(new_n802), .B2(new_n783), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1122), .A2(KEYINPUT125), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1107), .B1(new_n1122), .B2(KEYINPUT125), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(KEYINPUT126), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(KEYINPUT126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1120), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1106), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g704(.A1(G401), .A2(new_n462), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n655), .A2(new_n673), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g706(.A(new_n1132), .B1(new_n849), .B2(new_n851), .ZN(new_n1133));
  NAND2_X1  g707(.A1(new_n902), .A2(new_n1133), .ZN(G225));
  INV_X1    g708(.A(G225), .ZN(G308));
endmodule


