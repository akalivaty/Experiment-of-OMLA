//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  OR2_X1    g000(.A1(KEYINPUT69), .A2(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT69), .A2(G119), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G116), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(G116), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n192), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(new_n189), .C1(G116), .C2(new_n190), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT0), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT0), .B(G128), .Z(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(new_n198), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G137), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT66), .A4(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n206), .A2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT11), .B1(new_n204), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n212), .A2(new_n213), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n213), .B1(new_n212), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n203), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n198), .A2(G128), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI221_X1 g043(.A(KEYINPUT68), .B1(new_n224), .B2(new_n226), .C1(new_n198), .C2(G128), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n198), .A2(new_n224), .A3(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n216), .A2(new_n217), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n233), .A2(new_n234), .A3(G137), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n204), .B2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n205), .A2(new_n207), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(new_n215), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n212), .A2(new_n220), .A3(new_n213), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n223), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n197), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT70), .B(new_n203), .C1(new_n221), .C2(new_n222), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n246), .A2(KEYINPUT30), .A3(new_n241), .A4(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n246), .A2(new_n197), .A3(new_n241), .A4(new_n247), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n254), .B(new_n255), .Z(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT31), .B1(new_n249), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n242), .A2(new_n196), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n250), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n242), .A2(new_n196), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT28), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n259), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n250), .A2(new_n256), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n244), .A2(new_n248), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n258), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n258), .A2(new_n265), .A3(new_n270), .A4(KEYINPUT73), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(G472), .A2(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(KEYINPUT32), .A3(new_n276), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n262), .A2(new_n264), .A3(new_n259), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n267), .A2(new_n250), .ZN(new_n282));
  AOI211_X1 g096(.A(KEYINPUT29), .B(new_n281), .C1(new_n259), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n246), .A2(new_n241), .A3(new_n247), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n196), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n260), .B1(new_n285), .B2(new_n250), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(new_n264), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT29), .A3(new_n256), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G472), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n279), .A2(new_n280), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G140), .ZN(new_n294));
  INV_X1    g108(.A(G140), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G125), .ZN(new_n296));
  INV_X1    g110(.A(G146), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n295), .A2(KEYINPUT76), .A3(G125), .ZN(new_n301));
  XNOR2_X1  g115(.A(G125), .B(G140), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(KEYINPUT76), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n304));
  OAI211_X1 g118(.A(G146), .B(new_n300), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT69), .A2(G119), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT69), .A2(G119), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n308), .A2(new_n309), .A3(new_n200), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n187), .A2(G128), .A3(new_n188), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n200), .B1(new_n308), .B2(new_n309), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G110), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n200), .A2(G119), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n311), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n318), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT24), .B(G110), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n298), .B(new_n306), .C1(new_n321), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n316), .A2(new_n329), .A3(new_n320), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n317), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n294), .A2(new_n296), .A3(KEYINPUT76), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n295), .A2(KEYINPUT76), .A3(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  AOI21_X1  g149(.A(G146), .B1(new_n335), .B2(new_n300), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n306), .A2(new_n336), .B1(new_n322), .B2(new_n323), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n331), .A2(KEYINPUT77), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n316), .A2(new_n329), .A3(new_n320), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n329), .B1(new_n316), .B2(new_n320), .ZN(new_n341));
  OAI21_X1  g155(.A(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n337), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n326), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n346), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT77), .B1(new_n331), .B2(new_n337), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n343), .A3(new_n339), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n326), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n289), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G902), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n354), .B1(new_n353), .B2(new_n326), .ZN(new_n363));
  AOI211_X1 g177(.A(new_n325), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n362), .B(new_n289), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n358), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n362), .B1(new_n356), .B2(new_n289), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G214), .B1(G237), .B2(G902), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT82), .Z(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT83), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G122), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT8), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n189), .B(KEYINPUT5), .C1(G116), .C2(new_n190), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n375), .B(G113), .C1(KEYINPUT5), .C2(new_n189), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G107), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n380), .A2(G104), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n377), .A2(G107), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n376), .A2(new_n195), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n376), .B2(new_n195), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n374), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n347), .A2(G224), .ZN(new_n393));
  INV_X1    g207(.A(new_n231), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n228), .B2(new_n227), .ZN(new_n395));
  AOI21_X1  g209(.A(G125), .B1(new_n395), .B2(new_n230), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n203), .A2(G125), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT7), .B(new_n393), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n378), .A2(new_n381), .A3(new_n402), .A4(new_n383), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n382), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n196), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n389), .B(new_n373), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n232), .A2(new_n293), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n397), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n392), .A2(new_n399), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n289), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n389), .B1(new_n406), .B2(new_n408), .ZN(new_n415));
  INV_X1    g229(.A(new_n373), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n397), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n393), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n421), .A3(new_n416), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n414), .B1(new_n423), .B2(KEYINPUT84), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n418), .A2(new_n420), .A3(new_n425), .A4(new_n422), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n427), .B(KEYINPUT85), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n424), .B2(new_n426), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n372), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n212), .A2(new_n220), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n240), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n404), .A2(new_n407), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n203), .C1(new_n404), .C2(new_n405), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n388), .B1(new_n227), .B2(new_n394), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n384), .A2(new_n387), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n441), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n441), .A2(new_n442), .B1(new_n232), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n435), .A2(KEYINPUT80), .A3(new_n240), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n438), .A2(new_n440), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G140), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n347), .A2(G227), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n448), .B(new_n449), .Z(new_n450));
  AND2_X1   g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n229), .A2(new_n230), .A3(new_n231), .A4(new_n443), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n442), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT12), .B1(new_n436), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n435), .A2(new_n240), .B1(new_n452), .B2(new_n442), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(KEYINPUT12), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(KEYINPUT12), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n440), .A2(new_n445), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n436), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n447), .ZN(new_n464));
  INV_X1    g278(.A(new_n450), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n289), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n460), .A2(new_n447), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n465), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n451), .A2(new_n463), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(G469), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n468), .A2(new_n289), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT9), .B(G234), .ZN(new_n477));
  OAI21_X1  g291(.A(G221), .B1(new_n477), .B2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G113), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT90), .B(G104), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n334), .A2(new_n297), .B1(new_n298), .B2(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n303), .A2(G146), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(KEYINPUT87), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G214), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n486), .A2(G237), .A3(G953), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n487), .A2(G143), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT86), .B1(new_n487), .B2(G143), .ZN(new_n489));
  AND4_X1   g303(.A1(KEYINPUT86), .A2(new_n252), .A3(G143), .A4(G214), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT18), .A3(G131), .ZN(new_n492));
  AND2_X1   g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n485), .B(new_n492), .C1(new_n491), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(G131), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n488), .B(new_n213), .C1(new_n489), .C2(new_n490), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT19), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT19), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n302), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n297), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n305), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n305), .B2(new_n501), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n494), .B(KEYINPUT89), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n505), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n503), .A3(new_n497), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT89), .B1(new_n509), .B2(new_n494), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n482), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n306), .A2(new_n336), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n495), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n497), .A2(KEYINPUT17), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n494), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n482), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n511), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT20), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n511), .A2(new_n522), .A3(new_n518), .A4(new_n519), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n289), .B1(new_n516), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(G475), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n225), .A2(G128), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT13), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n225), .A3(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT92), .B1(new_n225), .B2(G128), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n200), .A3(G143), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n204), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n233), .A2(new_n537), .A3(new_n529), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT93), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n233), .A2(new_n537), .A3(new_n542), .A4(new_n529), .ZN(new_n543));
  XNOR2_X1  g357(.A(G116), .B(G122), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n380), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n539), .A2(new_n541), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT94), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n544), .B(G107), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n538), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n543), .A4(new_n541), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n537), .A2(new_n529), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n233), .ZN(new_n554));
  INV_X1    g368(.A(G122), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G116), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n380), .B1(new_n556), .B2(KEYINPUT14), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(new_n544), .Z(new_n558));
  NOR2_X1   g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n477), .A2(new_n357), .A3(G953), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n559), .B1(new_n547), .B2(new_n551), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n289), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n567), .B2(new_n289), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n347), .A2(G952), .ZN(new_n575));
  NAND2_X1  g389(.A1(G234), .A2(G237), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(G902), .A3(G953), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT21), .B(G898), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n524), .A2(new_n528), .A3(new_n574), .A4(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n433), .A2(new_n479), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n292), .A2(new_n369), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND2_X1  g401(.A1(new_n275), .A2(new_n289), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n589), .A2(new_n277), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n368), .A2(new_n479), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n567), .A2(new_n289), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT98), .B(G478), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT33), .B1(new_n565), .B2(KEYINPUT96), .ZN(new_n597));
  INV_X1    g411(.A(new_n566), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n565), .A2(new_n562), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n561), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n564), .A2(new_n602), .A3(KEYINPUT33), .A4(new_n566), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n568), .A2(G902), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n605), .A2(KEYINPUT97), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(KEYINPUT97), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n596), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n524), .A2(new_n528), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n583), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n371), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n427), .B1(new_n424), .B2(new_n426), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n428), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI211_X1 g428(.A(KEYINPUT95), .B(new_n427), .C1(new_n424), .C2(new_n426), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n593), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT99), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  AND2_X1   g435(.A1(new_n524), .A2(new_n528), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n572), .A2(new_n573), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n583), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n593), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  OR2_X1    g442(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n345), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n345), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n360), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n366), .B2(new_n367), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n585), .A2(new_n277), .A3(new_n589), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  INV_X1    g450(.A(new_n478), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n451), .A2(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(G902), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n474), .B1(new_n639), .B2(new_n468), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n637), .B1(new_n640), .B2(new_n473), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n641), .B(new_n611), .C1(new_n615), .C2(new_n614), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n623), .A2(new_n524), .A3(new_n528), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n577), .B(KEYINPUT100), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(new_n580), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n633), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n292), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT32), .B1(new_n275), .B2(new_n276), .ZN(new_n655));
  INV_X1    g469(.A(new_n276), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n278), .B(new_n656), .C1(new_n273), .C2(new_n274), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n650), .B1(new_n658), .B2(new_n291), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(KEYINPUT101), .A3(new_n643), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XNOR2_X1  g476(.A(new_n648), .B(KEYINPUT39), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n479), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT40), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n256), .B1(new_n285), .B2(new_n250), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n267), .B2(new_n266), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n667), .B2(G902), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n658), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n429), .A2(new_n432), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT38), .Z(new_n671));
  NOR4_X1   g485(.A1(new_n633), .A2(new_n622), .A3(new_n574), .A4(new_n371), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n665), .A2(new_n669), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  INV_X1    g488(.A(new_n633), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n658), .B2(new_n291), .ZN(new_n676));
  INV_X1    g490(.A(new_n648), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n608), .A2(new_n609), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n642), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(G469), .B1(new_n638), .B2(G902), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n469), .A2(new_n682), .A3(new_n478), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n292), .A2(new_n369), .A3(new_n617), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND4_X1  g501(.A1(new_n292), .A2(new_n369), .A3(new_n625), .A4(new_n684), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  INV_X1    g503(.A(new_n584), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n684), .B(new_n611), .C1(new_n614), .C2(new_n615), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n292), .A2(new_n690), .A3(new_n633), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  OAI211_X1 g508(.A(new_n258), .B(new_n270), .C1(new_n287), .C2(new_n256), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n588), .A2(G472), .B1(new_n276), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n574), .B1(new_n524), .B2(new_n528), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n611), .C1(new_n614), .C2(new_n615), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n683), .A2(new_n582), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n699), .A3(new_n369), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NAND2_X1  g516(.A1(new_n695), .A2(new_n276), .ZN(new_n703));
  AOI21_X1  g517(.A(G902), .B1(new_n273), .B2(new_n274), .ZN(new_n704));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n633), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n706), .A2(new_n678), .A3(new_n691), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n293), .ZN(G27));
  INV_X1    g522(.A(new_n678), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n469), .B(new_n475), .C1(new_n473), .C2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n710), .B2(new_n473), .ZN(new_n712));
  INV_X1    g526(.A(new_n432), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n428), .A3(new_n611), .A4(new_n478), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n292), .A2(new_n369), .A3(new_n709), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n279), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n655), .A2(KEYINPUT103), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n280), .A3(new_n291), .A4(new_n721), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n678), .A2(new_n712), .A3(new_n717), .A4(new_n714), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n369), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G131), .ZN(G33));
  NAND4_X1  g540(.A1(new_n292), .A2(new_n369), .A3(new_n649), .A4(new_n715), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  NAND2_X1  g542(.A1(new_n471), .A2(new_n472), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n733), .A3(G469), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n475), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n469), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT46), .B1(new_n735), .B2(new_n475), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n478), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(new_n663), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n608), .A2(new_n622), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n590), .A3(new_n675), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n670), .A2(new_n611), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT105), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n741), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n739), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT47), .B(new_n478), .C1(new_n737), .C2(new_n738), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n292), .A2(new_n369), .A3(new_n678), .A4(new_n749), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  NOR2_X1   g573(.A1(G952), .A2(G953), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n469), .A2(new_n682), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT106), .Z(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n637), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n755), .A3(new_n763), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n369), .A2(new_n744), .A3(new_n646), .A4(new_n696), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n750), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n714), .A2(new_n761), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n744), .A2(new_n767), .A3(new_n646), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n633), .A3(new_n696), .ZN(new_n769));
  INV_X1    g583(.A(new_n669), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(new_n369), .A3(new_n578), .A4(new_n767), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n608), .A2(new_n609), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n671), .A2(new_n611), .A3(new_n683), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n765), .A2(KEYINPUT50), .A3(new_n774), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n766), .A2(new_n779), .A3(KEYINPUT51), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n765), .A2(new_n692), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n608), .A2(new_n609), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n785), .B(new_n575), .C1(new_n786), .C2(new_n771), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n722), .A2(new_n369), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n768), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT48), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n768), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT110), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n787), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT48), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT110), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n784), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n787), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(KEYINPUT48), .A3(new_n790), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n784), .A2(new_n798), .A3(new_n799), .A4(new_n796), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n782), .B(new_n783), .C1(new_n797), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n707), .B1(new_n676), .B2(new_n679), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n648), .B(KEYINPUT108), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n712), .A2(new_n633), .A3(new_n637), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n669), .A2(new_n805), .A3(new_n699), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT101), .B1(new_n659), .B2(new_n643), .ZN(new_n807));
  AND4_X1   g621(.A1(KEYINPUT101), .A2(new_n292), .A3(new_n643), .A4(new_n651), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n803), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n661), .A2(KEYINPUT52), .A3(new_n806), .A4(new_n803), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n685), .A2(new_n688), .A3(new_n693), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n583), .B(new_n372), .C1(new_n429), .C2(new_n432), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n786), .B2(new_n644), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n277), .A3(new_n589), .A4(new_n591), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n586), .A2(new_n701), .A3(new_n817), .A4(new_n634), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n715), .A2(new_n696), .A3(new_n633), .A4(new_n709), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n479), .A2(new_n609), .A3(new_n623), .A4(new_n648), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n675), .A2(new_n749), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n292), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n727), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n725), .A2(new_n814), .A3(new_n818), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT107), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n685), .A2(new_n688), .A3(new_n693), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n586), .A2(new_n701), .A3(new_n817), .A4(new_n634), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT107), .A3(new_n725), .A4(new_n823), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n813), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n813), .A2(new_n826), .A3(KEYINPUT53), .A4(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n824), .A2(new_n832), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n831), .A2(new_n832), .B1(new_n813), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n838));
  AOI22_X1  g652(.A1(new_n835), .A2(KEYINPUT54), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n760), .B1(new_n802), .B2(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n762), .B(KEYINPUT49), .Z(new_n841));
  NAND4_X1  g655(.A1(new_n608), .A2(new_n622), .A3(new_n372), .A4(new_n478), .ZN(new_n842));
  OR4_X1    g656(.A1(new_n368), .A2(new_n841), .A3(new_n671), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n669), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT112), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  INV_X1    g660(.A(new_n844), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n837), .A2(new_n838), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n833), .B2(new_n834), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n801), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n846), .B(new_n847), .C1(new_n851), .C2(new_n760), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n852), .ZN(G75));
  NOR2_X1   g667(.A1(new_n347), .A2(G952), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n836), .A2(new_n813), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n833), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(G902), .A4(new_n430), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n418), .A2(new_n422), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(new_n420), .ZN(new_n861));
  XNOR2_X1  g675(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n864));
  NAND3_X1  g678(.A1(new_n859), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n837), .A2(new_n289), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n858), .B1(new_n866), .B2(new_n430), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n855), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n427), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n870), .A2(KEYINPUT114), .A3(new_n863), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT114), .B1(new_n870), .B2(new_n863), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G51));
  NOR2_X1   g687(.A1(new_n837), .A2(new_n838), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n848), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n475), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n467), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n837), .A2(new_n289), .A3(new_n735), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT118), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n854), .B1(new_n878), .B2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n511), .A2(new_n518), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n855), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(G60));
  AND2_X1   g699(.A1(new_n600), .A2(new_n603), .ZN(new_n886));
  NAND2_X1  g700(.A1(G478), .A2(G902), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n855), .B1(new_n875), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n839), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n891), .B2(new_n888), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(G63));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g708(.A1(G217), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT60), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  INV_X1    g712(.A(new_n896), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n837), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n356), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n855), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n630), .A2(new_n631), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n897), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n894), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n855), .A2(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n897), .A2(new_n900), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n904), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT120), .A4(new_n901), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n907), .A2(new_n914), .ZN(G66));
  INV_X1    g729(.A(G224), .ZN(new_n916));
  OAI21_X1  g730(.A(G953), .B1(new_n581), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n829), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n860), .B1(G898), .B2(new_n347), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n661), .A2(new_n803), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n788), .A2(new_n699), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n751), .B(new_n923), .C1(new_n740), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n758), .A2(new_n725), .A3(new_n727), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(G953), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n242), .A2(new_n243), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n248), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT122), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n498), .A2(new_n500), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(G900), .B2(G953), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n922), .B1(new_n927), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n347), .B1(G227), .B2(G900), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n923), .A2(new_n673), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n664), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n749), .B(new_n942), .C1(new_n786), .C2(new_n644), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n369), .A3(new_n292), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n941), .A2(new_n751), .A3(new_n758), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n933), .B1(new_n946), .B2(new_n347), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n937), .A2(new_n938), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n938), .B1(new_n937), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G72));
  XNOR2_X1  g764(.A(new_n282), .B(KEYINPUT127), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n256), .ZN(new_n952));
  INV_X1    g766(.A(new_n829), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n925), .A2(new_n953), .A3(new_n926), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n946), .A2(new_n953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(new_n957), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n256), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n958), .B(new_n855), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n282), .A2(new_n259), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n266), .A2(new_n267), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n835), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n962), .A2(new_n966), .ZN(G57));
endmodule


