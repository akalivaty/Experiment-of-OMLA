//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(G2104), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR3_X1   g038(.A1(new_n463), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(G101), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  OR2_X1    g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n467), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n463), .B2(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n460), .A2(new_n461), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n466), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n480), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n467), .A2(new_n469), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n479), .A2(new_n483), .ZN(G160));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n482), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n470), .A2(KEYINPUT69), .A3(new_n471), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT70), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  OAI221_X1 g069(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n482), .C2(G112), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n486), .A2(new_n461), .A3(new_n488), .ZN(new_n496));
  INV_X1    g071(.A(G136), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n494), .A2(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G114), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n503), .A3(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n509));
  OAI211_X1 g084(.A(G126), .B(G2105), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n482), .A2(new_n480), .A3(G138), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n482), .A2(new_n480), .A3(new_n514), .A4(G138), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(G164));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT72), .B1(new_n517), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(G651), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n522), .A2(G50), .A3(G543), .A4(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT5), .B(G543), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n520), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n519), .B1(KEYINPUT6), .B2(new_n520), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n517), .A2(KEYINPUT72), .A3(G651), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n527), .B(new_n523), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n518), .A2(new_n521), .B1(new_n517), .B2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n527), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n526), .B(new_n529), .C1(new_n530), .C2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  AND2_X1   g115(.A1(new_n536), .A2(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n527), .A2(G63), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n541), .A2(G51), .B1(G651), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n535), .A2(G89), .A3(new_n537), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G168));
  NAND3_X1  g123(.A1(new_n535), .A2(G90), .A3(new_n537), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n541), .A2(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT75), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n553), .A2(new_n554), .B1(G651), .B2(new_n556), .ZN(G171));
  AND2_X1   g132(.A1(new_n535), .A2(new_n537), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT5), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n541), .A2(G43), .B1(G651), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n535), .A2(G91), .A3(new_n537), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n527), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n520), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n522), .A2(G53), .A3(G543), .A4(new_n523), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT9), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n536), .A2(new_n582), .A3(G53), .A4(G543), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n581), .B1(new_n580), .B2(new_n583), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n576), .B(new_n578), .C1(new_n584), .C2(new_n585), .ZN(G299));
  NAND2_X1  g161(.A1(new_n553), .A2(new_n554), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n556), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G301));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n547), .B(new_n590), .ZN(G286));
  OAI21_X1  g166(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n536), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G49), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n558), .B2(G87), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G288));
  NAND4_X1  g172(.A1(new_n522), .A2(G48), .A3(G543), .A4(new_n523), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n536), .A2(KEYINPUT79), .A3(G48), .A4(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n535), .A2(G86), .A3(new_n537), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT78), .B1(new_n565), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n527), .A2(new_n607), .A3(G61), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n602), .A2(new_n603), .A3(new_n610), .ZN(G305));
  NAND2_X1  g186(.A1(new_n558), .A2(G85), .ZN(new_n612));
  NAND2_X1  g187(.A1(G72), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G60), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n565), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n541), .A2(G47), .B1(G651), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n558), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n538), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n619), .A2(new_n622), .B1(G54), .B2(new_n541), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G651), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n618), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n618), .B1(new_n627), .B2(G868), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(G868), .B2(new_n631), .ZN(G280));
  XOR2_X1   g207(.A(G280), .B(KEYINPUT81), .Z(G297));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n627), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g214(.A1(new_n482), .A2(G111), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n463), .B1(new_n640), .B2(KEYINPUT83), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n641), .B1(KEYINPUT83), .B2(new_n640), .C1(G99), .C2(G2105), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n493), .A2(G123), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n486), .A2(G135), .A3(new_n461), .A4(new_n488), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT84), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n476), .A2(new_n480), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT13), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XOR2_X1   g234(.A(G2427), .B(G2430), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT86), .B(KEYINPUT14), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  AND2_X1   g246(.A1(new_n671), .A2(G14), .ZN(G401));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT88), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT17), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n673), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(new_n676), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n673), .A3(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  INV_X1    g258(.A(new_n673), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n678), .A2(new_n684), .A3(new_n679), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n650), .ZN(new_n687));
  INV_X1    g262(.A(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n692), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n696), .A2(KEYINPUT20), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(new_n692), .A3(new_n695), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n699), .B(new_n701), .C1(KEYINPUT20), .C2(new_n696), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT89), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G5), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G171), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G1961), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  OAI221_X1 g292(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n482), .C2(G107), .ZN(new_n718));
  INV_X1    g293(.A(G131), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n496), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n493), .B2(G119), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n717), .B1(new_n721), .B2(new_n716), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G24), .ZN(new_n725));
  XNOR2_X1  g300(.A(G290), .B(KEYINPUT90), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(KEYINPUT36), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n711), .A2(G23), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n596), .B2(new_n711), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT92), .Z(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT33), .B(G1976), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n711), .A2(G22), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G166), .B2(new_n711), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G1971), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G1971), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n736), .A2(new_n737), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n711), .A2(G6), .ZN(new_n743));
  INV_X1    g318(.A(G305), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n711), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT32), .B(G1981), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT91), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT34), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT34), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n742), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n724), .B(new_n730), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(KEYINPUT93), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n749), .B(KEYINPUT34), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(KEYINPUT93), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n756), .A2(new_n757), .A3(new_n724), .A4(new_n730), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n716), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n716), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G2090), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n711), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n631), .B2(new_n711), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT102), .B(G1956), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT103), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT98), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT98), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n772), .A2(new_n487), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n486), .A2(G139), .A3(new_n461), .A4(new_n488), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n774), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n716), .ZN(new_n784));
  NOR2_X1   g359(.A1(G29), .A2(G33), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(KEYINPUT96), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT96), .B2(new_n785), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G2072), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G27), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G164), .B2(new_n716), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G2078), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT30), .B(G28), .Z(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT24), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n716), .B1(new_n794), .B2(G34), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(G34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G160), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n716), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n791), .B1(G29), .B2(new_n792), .C1(new_n793), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n711), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n569), .B2(new_n711), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n711), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n711), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n801), .A2(new_n793), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT31), .B(G11), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n806), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n649), .A2(new_n716), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n788), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n817));
  INV_X1    g392(.A(G140), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(new_n482), .B2(G116), .ZN(new_n819));
  NOR2_X1   g394(.A1(G104), .A2(G2105), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n496), .A2(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n493), .B2(G128), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n716), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n716), .A2(G26), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n817), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n817), .B2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(G2067), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n761), .A2(G2090), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n711), .A2(G4), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n627), .B2(new_n711), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT94), .B(G1348), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  AOI211_X1 g408(.A(new_n829), .B(new_n833), .C1(new_n828), .C2(new_n827), .ZN(new_n834));
  NOR2_X1   g409(.A1(G29), .A2(G32), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n476), .A2(G105), .ZN(new_n836));
  INV_X1    g411(.A(G141), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n496), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n493), .B2(G129), .ZN(new_n839));
  NAND3_X1  g414(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT26), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n835), .B1(new_n844), .B2(G29), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT27), .B(G1996), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND4_X1   g422(.A1(new_n770), .A2(new_n816), .A3(new_n834), .A4(new_n847), .ZN(new_n848));
  AND4_X1   g423(.A1(new_n715), .A2(new_n755), .A3(new_n758), .A4(new_n848), .ZN(G311));
  NAND4_X1  g424(.A1(new_n755), .A2(new_n758), .A3(new_n848), .A4(new_n715), .ZN(G150));
  NAND2_X1  g425(.A1(new_n558), .A2(G93), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n565), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n541), .A2(G55), .B1(G651), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n623), .A2(new_n626), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n634), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT39), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n856), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n569), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n858), .B1(new_n866), .B2(G860), .ZN(G145));
  OAI221_X1 g442(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n482), .C2(G118), .ZN(new_n868));
  INV_X1    g443(.A(G142), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n493), .A2(KEYINPUT106), .A3(G130), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n493), .B2(G130), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n868), .B1(new_n869), .B2(new_n496), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n721), .A2(new_n654), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n721), .A2(new_n654), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n844), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n843), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n513), .A2(new_n515), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n507), .A2(KEYINPUT105), .A3(new_n510), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  XNOR2_X1  g457(.A(KEYINPUT71), .B(G114), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n505), .B1(new_n883), .B2(G2105), .ZN(new_n884));
  INV_X1    g459(.A(new_n510), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n823), .B(new_n887), .Z(new_n888));
  AND3_X1   g463(.A1(new_n877), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n877), .B2(new_n879), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n873), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n877), .A2(new_n879), .ZN(new_n892));
  INV_X1    g467(.A(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n877), .A2(new_n879), .A3(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n872), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n783), .A2(G162), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n783), .A2(G162), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n897), .A2(new_n649), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n649), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n891), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n891), .B2(new_n896), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n800), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n891), .A2(new_n896), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(G160), .A3(new_n902), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n905), .A2(new_n909), .A3(new_n913), .A4(new_n910), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  NAND2_X1  g492(.A1(G303), .A2(new_n596), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(G303), .A2(new_n596), .ZN(new_n920));
  INV_X1    g495(.A(G290), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(G166), .A2(G288), .ZN(new_n923));
  AOI21_X1  g498(.A(G290), .B1(new_n923), .B2(new_n918), .ZN(new_n924));
  OAI21_X1  g499(.A(G305), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(G290), .A3(new_n918), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n744), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(new_n928), .ZN(new_n934));
  INV_X1    g509(.A(new_n931), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n932), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n569), .B(new_n856), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n636), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n627), .A2(G299), .ZN(new_n942));
  AOI21_X1  g517(.A(G299), .B1(new_n623), .B2(new_n626), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(KEYINPUT41), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n859), .A2(new_n631), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n947), .A2(new_n943), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(new_n941), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n938), .B1(new_n932), .B2(new_n936), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n939), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n939), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g532(.A(new_n956), .B1(G868), .B2(new_n864), .ZN(G331));
  NAND2_X1  g533(.A1(G286), .A2(G171), .ZN(new_n959));
  NAND2_X1  g534(.A1(G301), .A2(G168), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n940), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n940), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n951), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n960), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n865), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(new_n945), .A3(new_n948), .A4(new_n961), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n929), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n929), .A3(new_n967), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(KEYINPUT43), .A3(new_n910), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n910), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(KEYINPUT110), .A3(new_n910), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n976), .B2(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT44), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n969), .A2(new_n979), .A3(new_n910), .A4(new_n970), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n887), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(G40), .B1(new_n481), .B2(new_n482), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n477), .B1(new_n476), .B2(G101), .ZN(new_n990));
  INV_X1    g565(.A(G101), .ZN(new_n991));
  AOI211_X1 g566(.A(KEYINPUT68), .B(new_n991), .C1(new_n474), .C2(new_n475), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n473), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n823), .B(G2067), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n844), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n843), .A2(G1996), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n721), .A2(new_n723), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n721), .A2(new_n723), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1986), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(new_n921), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G290), .A2(G1986), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n995), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n479), .A2(new_n988), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G164), .B2(G1384), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n887), .B2(new_n985), .ZN(new_n1017));
  NOR3_X1   g592(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n994), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1019), .B2(G1956), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n580), .A2(new_n583), .ZN(new_n1023));
  AND4_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n576), .A4(new_n578), .ZN(new_n1024));
  AOI211_X1 g599(.A(new_n1021), .B(new_n1024), .C1(KEYINPUT57), .C2(G299), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1024), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT115), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1020), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1024), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n1015), .C1(new_n1019), .C2(G1956), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(KEYINPUT61), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1033));
  INV_X1    g608(.A(new_n1031), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n514), .B1(new_n472), .B2(G138), .ZN(new_n1035));
  INV_X1    g610(.A(new_n515), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n507), .B(new_n510), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1016), .A3(new_n985), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n507), .A2(KEYINPUT105), .A3(new_n510), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT105), .B1(new_n507), .B2(new_n510), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1384), .B1(new_n1041), .B2(new_n880), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1011), .B(new_n1038), .C1(new_n1042), .C2(new_n1016), .ZN(new_n1043));
  INV_X1    g618(.A(G1956), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1030), .B1(new_n1045), .B2(new_n1015), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1033), .B1(new_n1034), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n985), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n994), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n886), .A2(new_n881), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1016), .B(new_n985), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n887), .A2(KEYINPUT111), .A3(new_n1016), .A4(new_n985), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1011), .A2(new_n887), .A3(new_n985), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1056), .A2(new_n832), .B1(new_n828), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n627), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1032), .A2(new_n1047), .A3(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1010), .A2(new_n998), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n1063), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n569), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1072), .A3(new_n569), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT59), .A3(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1069), .A2(new_n569), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT119), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1071), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n1073), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1059), .A2(new_n859), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1059), .A2(new_n859), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT60), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1062), .A2(new_n1078), .A3(new_n1079), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1029), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1031), .B1(new_n1084), .B2(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT116), .B(new_n1031), .C1(new_n1084), .C2(new_n1081), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT122), .B1(new_n993), .B2(new_n473), .ZN(new_n1091));
  AND4_X1   g666(.A1(KEYINPUT122), .A2(new_n466), .A3(new_n473), .A4(new_n478), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n989), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT123), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(new_n989), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n987), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT124), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G2078), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1094), .A2(new_n1101), .A3(new_n987), .A4(new_n1096), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1098), .A2(new_n1010), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1056), .A2(new_n714), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1099), .B1(new_n1105), .B2(G2078), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(G301), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n986), .B2(new_n994), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT113), .B(new_n1011), .C1(new_n1042), .C2(KEYINPUT45), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1037), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1100), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1104), .B(new_n1106), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1108), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT125), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1120), .B(KEYINPUT54), .C1(new_n1108), .C2(new_n1116), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1113), .A2(new_n809), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(KEYINPUT114), .A3(new_n793), .A4(new_n1049), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1056), .B2(G2084), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G8), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n547), .A2(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1128), .A2(G8), .A3(new_n547), .ZN(new_n1135));
  OAI211_X1 g710(.A(G8), .B(new_n1132), .C1(new_n1128), .C2(new_n547), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1971), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1105), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1056), .B2(G2090), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(G8), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G303), .A2(G8), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT55), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G2090), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1019), .A2(new_n1145), .B1(new_n1138), .B2(new_n1105), .ZN(new_n1146));
  INV_X1    g721(.A(G8), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(G305), .A2(G1981), .ZN(new_n1149));
  INV_X1    g724(.A(G1981), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n602), .A2(new_n603), .A3(new_n610), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT49), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1058), .A2(new_n1147), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1149), .A2(KEYINPUT49), .A3(new_n1151), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1976), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT52), .B1(G288), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n596), .A2(G1976), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(G8), .A3(new_n1057), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT52), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT112), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1144), .B(new_n1148), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1103), .A2(KEYINPUT126), .A3(new_n1107), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(G171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1115), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1118), .B1(new_n1174), .B2(G301), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1168), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1090), .A2(new_n1122), .A3(new_n1137), .A4(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(new_n1164), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1129), .A2(G286), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT63), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1144), .A2(new_n1164), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1157), .A2(new_n1158), .A3(new_n596), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1151), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1155), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1177), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1116), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1134), .A2(new_n1190), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1180), .A2(KEYINPUT63), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1168), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1009), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n995), .A2(new_n998), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT46), .Z(new_n1197));
  NAND2_X1  g772(.A1(new_n996), .A2(new_n844), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n995), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT47), .Z(new_n1200));
  NOR4_X1   g775(.A1(new_n997), .A2(new_n999), .A3(new_n1003), .A4(new_n1000), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n823), .A2(new_n828), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n995), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1004), .A2(new_n995), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n995), .A2(new_n1008), .ZN(new_n1206));
  XOR2_X1   g781(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1207));
  XNOR2_X1  g782(.A(new_n1206), .B(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1204), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1195), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(G319), .ZN(new_n1212));
  NOR2_X1   g786(.A1(G401), .A2(new_n1212), .ZN(new_n1213));
  AND3_X1   g787(.A1(new_n689), .A2(new_n911), .A3(new_n1213), .ZN(new_n1214));
  AND3_X1   g788(.A1(new_n1214), .A2(new_n709), .A3(new_n981), .ZN(G308));
  NAND3_X1  g789(.A1(new_n1214), .A2(new_n981), .A3(new_n709), .ZN(G225));
endmodule


