//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n452), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(new_n463), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n478), .ZN(G160));
  AOI21_X1  g054(.A(new_n472), .B1(new_n464), .B2(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n472), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(G136), .B2(new_n467), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(G162));
  NOR2_X1   g061(.A1(new_n472), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n480), .B2(G126), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n467), .B2(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n491), .A2(G138), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT70), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n503), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n503), .A2(G543), .A3(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(new_n498), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n511), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n503), .A2(G543), .A3(new_n510), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n509), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n520), .A2(new_n522), .A3(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n509), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n511), .A2(new_n534), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n537), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n533), .B1(new_n539), .B2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n519), .A2(G81), .B1(new_n521), .B2(G43), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n498), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  AND2_X1   g127(.A1(new_n519), .A2(G91), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(G543), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n506), .A2(new_n558), .A3(new_n508), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n554), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(G78), .A2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n564), .B(G651), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n553), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n503), .A2(G53), .A3(G543), .A4(new_n510), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT73), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n521), .A2(new_n574), .A3(new_n575), .A4(G53), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n499), .A2(new_n502), .B1(KEYINPUT6), .B2(new_n498), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n577), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n572), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n573), .B1(new_n572), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n566), .B1(new_n581), .B2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n519), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n521), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n498), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n519), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n521), .A2(G48), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n511), .A2(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n498), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(G290));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n511), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n577), .A2(KEYINPUT10), .A3(G92), .A4(new_n509), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n557), .B2(new_n559), .ZN(new_n610));
  AND2_X1   g185(.A1(G79), .A2(G543), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n513), .A2(KEYINPUT79), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n577), .A2(new_n614), .A3(G543), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(G54), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n608), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT80), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n608), .A2(new_n612), .A3(new_n619), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  MUX2_X1   g198(.A(G301), .B(new_n622), .S(new_n623), .Z(G284));
  MUX2_X1   g199(.A(G301), .B(new_n622), .S(new_n623), .Z(G321));
  NAND2_X1  g200(.A1(G299), .A2(new_n623), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n623), .B2(G168), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(new_n623), .B2(G168), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n621), .B1(new_n629), .B2(G860), .ZN(G148));
  AOI21_X1  g205(.A(KEYINPUT81), .B1(new_n621), .B2(new_n629), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n632));
  AOI211_X1 g207(.A(new_n632), .B(G559), .C1(new_n618), .C2(new_n620), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n631), .A2(new_n633), .A3(new_n623), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n623), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n493), .A2(G2104), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n467), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n480), .A2(G123), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT82), .Z(G156));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n656), .A2(KEYINPUT85), .A3(KEYINPUT14), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT85), .B1(new_n656), .B2(KEYINPUT14), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n660), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n655), .B(new_n665), .C1(new_n657), .C2(new_n658), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n661), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n661), .B2(new_n666), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n650), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n670), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(new_n668), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(KEYINPUT86), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(KEYINPUT86), .B2(new_n676), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n675), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n676), .B(new_n682), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n678), .B(new_n680), .C1(new_n681), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n679), .A2(new_n676), .A3(new_n675), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(new_n681), .A3(new_n679), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  XOR2_X1   g275(.A(G1961), .B(G1966), .Z(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(new_n703), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n699), .A2(new_n702), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n709), .B1(new_n706), .B2(new_n708), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n696), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(new_n696), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n714), .A2(new_n715), .A3(new_n710), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n713), .B2(new_n716), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(G229));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G24), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  INV_X1    g300(.A(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n480), .A2(G119), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G107), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n467), .B2(G131), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XOR2_X1   g315(.A(new_n739), .B(new_n740), .Z(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G23), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT92), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G288), .B2(new_n721), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT33), .B(G1976), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n721), .A2(G22), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G166), .B2(new_n721), .ZN(new_n750));
  INV_X1    g325(.A(G1971), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G6), .B(G305), .S(G16), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT32), .B(G1981), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n747), .A2(new_n748), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n727), .B(new_n741), .C1(new_n756), .C2(KEYINPUT34), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(KEYINPUT34), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n757), .A2(new_n758), .B1(KEYINPUT94), .B2(KEYINPUT36), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT95), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n721), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1956), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n621), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1348), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G35), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G162), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(G160), .A2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n776), .B2(KEYINPUT24), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(KEYINPUT24), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n728), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n467), .A2(G141), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT26), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(G105), .B2(new_n469), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n480), .A2(G129), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n781), .B1(new_n792), .B2(new_n728), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT98), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n780), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n728), .A2(G33), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT25), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n467), .A2(G139), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(new_n472), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n797), .B1(new_n804), .B2(new_n728), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G2072), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(G2072), .ZN(new_n807));
  INV_X1    g382(.A(G28), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT30), .ZN(new_n809));
  AOI21_X1  g384(.A(G29), .B1(new_n808), .B2(KEYINPUT30), .ZN(new_n810));
  OR2_X1    g385(.A1(KEYINPUT31), .A2(G11), .ZN(new_n811));
  NAND2_X1  g386(.A1(KEYINPUT31), .A2(G11), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n807), .B(new_n813), .C1(new_n728), .C2(new_n646), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n796), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n721), .A2(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n547), .B2(new_n721), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1341), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n728), .A2(G26), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT28), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n480), .A2(G128), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n472), .A2(G116), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n467), .A2(G140), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT96), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n467), .A2(new_n827), .A3(G140), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n824), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n820), .B1(new_n830), .B2(G29), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2067), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n774), .A2(new_n815), .A3(new_n818), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G168), .A2(G16), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G21), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(KEYINPUT99), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(KEYINPUT99), .B2(new_n834), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1966), .ZN(new_n838));
  NOR2_X1   g413(.A1(G164), .A2(new_n728), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G27), .B2(new_n728), .ZN(new_n840));
  INV_X1    g415(.A(G2078), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n793), .A2(new_n795), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n838), .B(new_n842), .C1(new_n841), .C2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n721), .A2(G5), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G171), .B2(new_n721), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1961), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n773), .A2(G2090), .ZN(new_n847));
  NOR4_X1   g422(.A1(new_n833), .A2(new_n843), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n762), .A2(new_n766), .A3(new_n770), .A4(new_n848), .ZN(G150));
  INV_X1    g424(.A(G150), .ZN(G311));
  AOI22_X1  g425(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT101), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(G651), .A3(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n519), .A2(G93), .B1(new_n521), .B2(G55), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n621), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n854), .A2(new_n545), .A3(new_n543), .A4(new_n855), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n854), .A2(new_n855), .B1(new_n543), .B2(new_n545), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n861), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT102), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n866), .B2(new_n867), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n858), .B1(new_n869), .B2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(G160), .B(new_n646), .ZN(new_n873));
  XNOR2_X1  g448(.A(G162), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n738), .B(new_n638), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n467), .A2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n480), .A2(G130), .ZN(new_n878));
  OR2_X1    g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n804), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n496), .A2(KEYINPUT103), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(new_n490), .C1(new_n492), .C2(new_n495), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n829), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n829), .B1(new_n885), .B2(new_n887), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n889), .A2(new_n890), .A3(new_n791), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n830), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n792), .B1(new_n893), .B2(new_n888), .ZN(new_n894));
  OAI211_X1 g469(.A(KEYINPUT104), .B(new_n884), .C1(new_n891), .C2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n791), .B1(new_n889), .B2(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n792), .A3(new_n888), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n883), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n883), .B1(new_n895), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n875), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n895), .A2(new_n900), .ZN(new_n905));
  INV_X1    g480(.A(new_n883), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n883), .A2(new_n895), .A3(new_n900), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n874), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g486(.A(KEYINPUT108), .B1(new_n856), .B2(new_n623), .ZN(new_n912));
  INV_X1    g487(.A(new_n865), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n631), .B2(new_n633), .ZN(new_n914));
  INV_X1    g489(.A(G54), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n513), .B2(KEYINPUT79), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n606), .A2(new_n607), .B1(new_n916), .B2(new_n615), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n619), .B1(new_n917), .B2(new_n612), .ZN(new_n918));
  INV_X1    g493(.A(new_n620), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n629), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n632), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n621), .A2(KEYINPUT81), .A3(new_n629), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n865), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n914), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n617), .ZN(new_n925));
  NAND2_X1  g500(.A1(G299), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n566), .B(new_n617), .C1(new_n581), .C2(new_n582), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(KEYINPUT105), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT105), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT9), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n570), .B1(new_n567), .B2(KEYINPUT9), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT75), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n572), .A2(new_n580), .A3(new_n573), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n941), .A2(KEYINPUT106), .A3(new_n566), .A4(new_n617), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n933), .A2(new_n926), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(G299), .B2(new_n925), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n927), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n931), .B1(new_n924), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(G290), .B(G305), .ZN(new_n948));
  XOR2_X1   g523(.A(G166), .B(G288), .Z(new_n949));
  OR2_X1    g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n949), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n931), .B(new_n953), .C1(new_n924), .C2(new_n946), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G868), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n955), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n912), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(KEYINPUT108), .A3(G868), .A4(new_n959), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(G295));
  AND2_X1   g540(.A1(new_n962), .A2(new_n964), .ZN(G331));
  NAND2_X1  g541(.A1(new_n856), .A2(new_n546), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n967), .A2(G301), .A3(new_n862), .ZN(new_n968));
  AOI21_X1  g543(.A(G301), .B1(new_n967), .B2(new_n862), .ZN(new_n969));
  OAI21_X1  g544(.A(G286), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(G171), .B1(new_n863), .B2(new_n864), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(G301), .A3(new_n862), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(G168), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n926), .A2(new_n927), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n946), .B2(new_n974), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n948), .B(new_n949), .Z(new_n978));
  AOI21_X1  g553(.A(G37), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n950), .A2(new_n952), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n976), .C1(new_n946), .C2(new_n974), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT43), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n928), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n983), .B2(new_n929), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(new_n944), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n945), .A2(new_n933), .A3(new_n942), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n973), .A4(new_n970), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n978), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n981), .A3(new_n904), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT44), .B1(new_n982), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n979), .B2(new_n981), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n988), .A2(new_n981), .A3(new_n990), .A4(new_n904), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n996), .B2(KEYINPUT44), .ZN(G397));
  OAI21_X1  g572(.A(KEYINPUT109), .B1(new_n892), .B2(G1384), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n885), .A2(new_n1000), .A3(new_n1001), .A4(new_n887), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n478), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(G40), .A3(new_n468), .A4(new_n470), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n791), .B(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n829), .B(G2067), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n738), .B(new_n740), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n496), .A2(new_n1001), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1005), .B1(new_n1015), .B2(new_n999), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n1001), .A4(new_n887), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n496), .A2(KEYINPUT110), .A3(new_n1001), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT110), .B1(new_n496), .B2(new_n1001), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1005), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n496), .A2(new_n1027), .A3(new_n1001), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT113), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n496), .A2(new_n1030), .A3(new_n1027), .A4(new_n1001), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1026), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1956), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1019), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT57), .B1(new_n572), .B2(new_n580), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n566), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1035), .A2(KEYINPUT118), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1035), .A2(KEYINPUT118), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1015), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n1022), .A3(new_n1020), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1005), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1348), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1026), .A3(new_n1022), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2067), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n621), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1052), .B(KEYINPUT117), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1040), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1016), .A2(new_n1017), .A3(new_n1007), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1056), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1055), .B(new_n547), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1061), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(new_n1059), .A3(new_n1058), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(KEYINPUT121), .A3(new_n1055), .A4(new_n547), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n547), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(KEYINPUT59), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1069), .B2(KEYINPUT59), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1039), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1049), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1051), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1082), .A2(new_n1083), .B1(KEYINPUT60), .B2(new_n621), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1076), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1054), .B1(new_n1073), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G86), .ZN(new_n1087));
  INV_X1    g662(.A(G48), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n511), .A2(new_n1087), .B1(new_n513), .B2(new_n1088), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n1089), .A2(new_n591), .A3(G1981), .ZN(new_n1090));
  OAI21_X1  g665(.A(G1981), .B1(new_n1089), .B2(new_n591), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(KEYINPUT49), .A3(new_n1091), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(G8), .A3(new_n1050), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G288), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G1976), .ZN(new_n1098));
  INV_X1    g673(.A(G1976), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1050), .A2(G8), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1050), .A2(G8), .A3(new_n1098), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(KEYINPUT52), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n751), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(G2090), .ZN(new_n1108));
  INV_X1    g683(.A(G8), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G166), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT55), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT112), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1113), .A3(KEYINPUT55), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(new_n1114), .C1(KEYINPUT55), .C2(new_n1110), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1108), .A2(new_n1115), .A3(G8), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1104), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1106), .B1(new_n1033), .B2(G2090), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(G8), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1961), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1107), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1016), .A2(new_n1017), .A3(new_n841), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  AOI21_X1  g699(.A(G171), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n999), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1126));
  OAI211_X1 g701(.A(G40), .B(G160), .C1(new_n1015), .C2(new_n999), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .A4(new_n841), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT53), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1046), .A2(new_n1022), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1132), .B2(new_n999), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n1133), .B2(new_n841), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1122), .B(new_n1125), .C1(new_n1131), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT124), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1005), .A2(new_n1124), .A3(G2078), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1003), .A2(new_n1017), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n1122), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1141), .B2(G171), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1126), .A2(new_n1128), .A3(new_n841), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT53), .A3(new_n1130), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1136), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1966), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT45), .B1(new_n1046), .B2(new_n1022), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1127), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT114), .B(G2084), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1047), .A2(new_n1048), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(G168), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G8), .ZN(new_n1155));
  AOI21_X1  g730(.A(G168), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT51), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(KEYINPUT51), .B2(new_n1155), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1120), .A2(new_n1148), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1140), .B(new_n1122), .C1(new_n1131), .C2(new_n1134), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(G171), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1139), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1137), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1086), .A2(new_n1159), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(KEYINPUT62), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1157), .B(new_n1171), .C1(KEYINPUT51), .C2(new_n1155), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n1120), .A4(new_n1172), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1109), .B(G286), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1108), .A2(G8), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT63), .B(new_n1174), .C1(new_n1175), .C2(new_n1115), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT116), .B1(new_n1176), .B2(new_n1117), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1115), .B1(new_n1108), .B2(G8), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(G8), .A3(G168), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT116), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n1116), .A4(new_n1104), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1117), .A2(new_n1119), .A3(new_n1180), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1177), .B(new_n1184), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1050), .A2(G8), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1096), .A2(new_n1099), .A3(new_n1097), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n1189), .B2(new_n1090), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1116), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1191), .B2(new_n1104), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1173), .A2(new_n1187), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1014), .B1(new_n1168), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT46), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1009), .B(new_n792), .C1(new_n1195), .C2(G1996), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1006), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1198), .A2(KEYINPUT125), .A3(new_n1195), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT125), .B1(new_n1198), .B2(new_n1195), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT47), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1006), .A2(new_n726), .A3(new_n724), .ZN(new_n1205));
  XNOR2_X1  g780(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1006), .A2(new_n1012), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1010), .A2(new_n740), .A3(new_n733), .A4(new_n737), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(G2067), .B2(new_n830), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1207), .A2(new_n1208), .B1(new_n1210), .B2(new_n1006), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1203), .A2(new_n1204), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1194), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n943), .A2(new_n944), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n945), .A2(new_n927), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n974), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g792(.A1(new_n974), .A2(new_n975), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n978), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1220), .A2(new_n904), .A3(new_n981), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1221), .A2(KEYINPUT43), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1222), .A2(new_n994), .ZN(new_n1223));
  NOR2_X1   g797(.A1(G227), .A2(new_n460), .ZN(new_n1224));
  OAI21_X1  g798(.A(new_n1224), .B1(new_n718), .B2(new_n719), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1225), .B1(new_n671), .B2(new_n673), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n910), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g801(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1215), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g803(.A(KEYINPUT127), .B(new_n1227), .C1(new_n1222), .C2(new_n994), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1229), .A2(new_n1230), .ZN(G308));
  OAI21_X1  g805(.A(KEYINPUT127), .B1(new_n996), .B2(new_n1227), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1223), .A2(new_n1215), .A3(new_n1228), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1233), .ZN(G225));
endmodule


