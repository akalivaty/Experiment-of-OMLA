

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XNOR2_X2 U326 ( .A(n406), .B(n405), .ZN(n557) );
  XNOR2_X1 U327 ( .A(n294), .B(KEYINPUT55), .ZN(n460) );
  AND2_X1 U328 ( .A1(n576), .A2(n476), .ZN(n294) );
  INV_X1 U329 ( .A(KEYINPUT54), .ZN(n424) );
  XNOR2_X1 U330 ( .A(n295), .B(n363), .ZN(n370) );
  XNOR2_X1 U331 ( .A(n383), .B(n382), .ZN(n387) );
  INV_X1 U332 ( .A(KEYINPUT48), .ZN(n405) );
  XOR2_X1 U333 ( .A(n390), .B(KEYINPUT31), .Z(n295) );
  XOR2_X1 U334 ( .A(n448), .B(n378), .Z(n296) );
  XOR2_X1 U335 ( .A(n367), .B(n366), .Z(n297) );
  INV_X1 U336 ( .A(KEYINPUT9), .ZN(n380) );
  XNOR2_X1 U337 ( .A(n368), .B(n297), .ZN(n369) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G106GAT), .ZN(n361) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U340 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U341 ( .A(n362), .B(n361), .ZN(n390) );
  XOR2_X1 U342 ( .A(n372), .B(n371), .Z(n583) );
  XOR2_X1 U343 ( .A(KEYINPUT77), .B(n570), .Z(n551) );
  NOR2_X2 U344 ( .A1(n460), .A2(n472), .ZN(n573) );
  XNOR2_X1 U345 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U346 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U347 ( .A(G57GAT), .B(KEYINPUT88), .Z(n299) );
  XNOR2_X1 U348 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U350 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n301) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(KEYINPUT87), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U353 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U354 ( .A(KEYINPUT0), .B(G127GAT), .Z(n450) );
  XOR2_X1 U355 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n305) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n450), .B(n306), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U360 ( .A(G85GAT), .B(G162GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U363 ( .A(n312), .B(n311), .Z(n321) );
  XOR2_X1 U364 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n314) );
  XNOR2_X1 U365 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(n315), .ZN(n443) );
  INV_X1 U368 ( .A(n443), .ZN(n319) );
  XOR2_X1 U369 ( .A(KEYINPUT1), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G120GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n528) );
  XOR2_X1 U374 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n323) );
  XNOR2_X1 U375 ( .A(KEYINPUT14), .B(KEYINPUT79), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n331) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n329) );
  XOR2_X1 U378 ( .A(G78GAT), .B(G211GAT), .Z(n325) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G127GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U381 ( .A(G183GAT), .B(G71GAT), .Z(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n339) );
  XNOR2_X1 U385 ( .A(G22GAT), .B(G1GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n332), .B(G8GAT), .ZN(n346) );
  XOR2_X1 U387 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n334) );
  XNOR2_X1 U388 ( .A(G155GAT), .B(G64GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n346), .B(n335), .ZN(n337) );
  XOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT13), .Z(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT69), .B(n336), .Z(n354) );
  XOR2_X1 U393 ( .A(n337), .B(n354), .Z(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n587) );
  XOR2_X1 U395 ( .A(G141GAT), .B(G197GAT), .Z(n341) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(G50GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n353) );
  XOR2_X1 U398 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n343) );
  NAND2_X1 U399 ( .A1(G229GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U401 ( .A(n344), .B(KEYINPUT29), .Z(n348) );
  XNOR2_X1 U402 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n345), .B(KEYINPUT7), .ZN(n378) );
  XNOR2_X1 U404 ( .A(n378), .B(n346), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U406 ( .A(G113GAT), .B(G15GAT), .Z(n451) );
  XOR2_X1 U407 ( .A(n349), .B(n451), .Z(n351) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G43GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U410 ( .A(n353), .B(n352), .Z(n577) );
  INV_X1 U411 ( .A(n577), .ZN(n560) );
  XOR2_X1 U412 ( .A(n354), .B(G92GAT), .Z(n356) );
  XOR2_X1 U413 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XNOR2_X1 U414 ( .A(G176GAT), .B(n445), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n372) );
  INV_X1 U416 ( .A(G85GAT), .ZN(n357) );
  NAND2_X1 U417 ( .A1(n357), .A2(KEYINPUT73), .ZN(n360) );
  INV_X1 U418 ( .A(KEYINPUT73), .ZN(n358) );
  NAND2_X1 U419 ( .A1(n358), .A2(G85GAT), .ZN(n359) );
  NAND2_X1 U420 ( .A1(n360), .A2(n359), .ZN(n362) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n364), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U424 ( .A(G204GAT), .B(G64GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n365), .B(KEYINPUT74), .ZN(n413) );
  XNOR2_X1 U426 ( .A(n439), .B(n413), .ZN(n368) );
  XOR2_X1 U427 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n367) );
  XNOR2_X1 U428 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n583), .B(KEYINPUT64), .ZN(n374) );
  INV_X1 U430 ( .A(KEYINPUT41), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n563) );
  AND2_X1 U432 ( .A1(n560), .A2(n563), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n375), .B(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U434 ( .A1(n587), .A2(n376), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n377), .B(KEYINPUT113), .ZN(n393) );
  XOR2_X1 U436 ( .A(G43GAT), .B(G134GAT), .Z(n448) );
  NAND2_X1 U437 ( .A1(G232GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n296), .B(n379), .ZN(n383) );
  XOR2_X1 U439 ( .A(G50GAT), .B(G162GAT), .Z(n432) );
  XNOR2_X1 U440 ( .A(n432), .B(KEYINPUT10), .ZN(n381) );
  XOR2_X1 U441 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT66), .B(KEYINPUT75), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U445 ( .A(G92GAT), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(G190GAT), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n410) );
  XOR2_X1 U448 ( .A(n390), .B(n410), .Z(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n570) );
  NOR2_X1 U450 ( .A1(n393), .A2(n570), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(KEYINPUT47), .ZN(n404) );
  XNOR2_X1 U452 ( .A(n551), .B(KEYINPUT103), .ZN(n395) );
  NAND2_X1 U453 ( .A1(n395), .A2(KEYINPUT36), .ZN(n399) );
  INV_X1 U454 ( .A(n395), .ZN(n397) );
  INV_X1 U455 ( .A(KEYINPUT36), .ZN(n396) );
  NAND2_X1 U456 ( .A1(n397), .A2(n396), .ZN(n398) );
  NAND2_X1 U457 ( .A1(n399), .A2(n398), .ZN(n498) );
  INV_X1 U458 ( .A(n587), .ZN(n500) );
  NOR2_X1 U459 ( .A1(n498), .A2(n500), .ZN(n400) );
  XOR2_X1 U460 ( .A(n400), .B(KEYINPUT45), .Z(n401) );
  NOR2_X1 U461 ( .A1(n583), .A2(n401), .ZN(n402) );
  NAND2_X1 U462 ( .A1(n402), .A2(n577), .ZN(n403) );
  NAND2_X1 U463 ( .A1(n404), .A2(n403), .ZN(n406) );
  XOR2_X1 U464 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n408) );
  NAND2_X1 U465 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U467 ( .A(KEYINPUT93), .B(n409), .Z(n412) );
  XNOR2_X1 U468 ( .A(G8GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n422) );
  XOR2_X1 U471 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n416) );
  XNOR2_X1 U472 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U474 ( .A(n417), .B(G183GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(G176GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n457) );
  XNOR2_X1 U477 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n420), .B(G211GAT), .ZN(n440) );
  XNOR2_X1 U479 ( .A(n457), .B(n440), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n531) );
  XNOR2_X1 U481 ( .A(KEYINPUT121), .B(n531), .ZN(n423) );
  NOR2_X1 U482 ( .A1(n557), .A2(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U484 ( .A1(n528), .A2(n426), .ZN(n428) );
  INV_X1 U485 ( .A(KEYINPUT65), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n576) );
  XOR2_X1 U487 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n430) );
  XNOR2_X1 U488 ( .A(G218GAT), .B(G106GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT86), .B(G204GAT), .Z(n436) );
  XNOR2_X1 U494 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U496 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n476) );
  XOR2_X1 U500 ( .A(n445), .B(KEYINPUT83), .Z(n447) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n453) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n459) );
  XOR2_X1 U506 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n455) );
  XNOR2_X1 U507 ( .A(G190GAT), .B(G99GAT), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U509 ( .A(n457), .B(n456), .Z(n458) );
  XNOR2_X1 U510 ( .A(n459), .B(n458), .ZN(n472) );
  NAND2_X1 U511 ( .A1(n573), .A2(n563), .ZN(n463) );
  XOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U514 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NAND2_X1 U515 ( .A1(n560), .A2(n573), .ZN(n465) );
  XNOR2_X1 U516 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n465), .B(n464), .ZN(G1348GAT) );
  NAND2_X1 U518 ( .A1(n573), .A2(n551), .ZN(n468) );
  XOR2_X1 U519 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT84), .B(n472), .ZN(n470) );
  XNOR2_X1 U521 ( .A(n476), .B(KEYINPUT67), .ZN(n469) );
  XNOR2_X1 U522 ( .A(n469), .B(KEYINPUT28), .ZN(n537) );
  XNOR2_X1 U523 ( .A(n531), .B(KEYINPUT27), .ZN(n478) );
  NAND2_X1 U524 ( .A1(n528), .A2(n478), .ZN(n556) );
  NOR2_X1 U525 ( .A1(n537), .A2(n556), .ZN(n541) );
  NAND2_X1 U526 ( .A1(n470), .A2(n541), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n471), .B(KEYINPUT95), .ZN(n484) );
  INV_X1 U528 ( .A(n472), .ZN(n542) );
  AND2_X1 U529 ( .A1(n531), .A2(n542), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(n473), .Z(n474) );
  NAND2_X1 U531 ( .A1(n476), .A2(n474), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(n475), .Z(n480) );
  NOR2_X1 U533 ( .A1(n542), .A2(n476), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT26), .B(n477), .ZN(n575) );
  NAND2_X1 U535 ( .A1(n478), .A2(n575), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT97), .B(n481), .ZN(n482) );
  NOR2_X1 U538 ( .A1(n482), .A2(n528), .ZN(n483) );
  NOR2_X1 U539 ( .A1(n484), .A2(n483), .ZN(n499) );
  NOR2_X1 U540 ( .A1(n551), .A2(n500), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(n485), .Z(n486) );
  NOR2_X1 U542 ( .A1(n499), .A2(n486), .ZN(n487) );
  XOR2_X1 U543 ( .A(KEYINPUT98), .B(n487), .Z(n515) );
  OR2_X1 U544 ( .A1(n577), .A2(n583), .ZN(n503) );
  NOR2_X1 U545 ( .A1(n515), .A2(n503), .ZN(n496) );
  NAND2_X1 U546 ( .A1(n496), .A2(n528), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n489) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  XOR2_X1 U551 ( .A(G8GAT), .B(KEYINPUT101), .Z(n493) );
  NAND2_X1 U552 ( .A1(n496), .A2(n531), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U555 ( .A1(n496), .A2(n542), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n496), .A2(n537), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n506) );
  NOR2_X1 U560 ( .A1(n498), .A2(n499), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U562 ( .A(KEYINPUT37), .B(n502), .Z(n527) );
  OR2_X1 U563 ( .A1(n527), .A2(n503), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT38), .B(n504), .Z(n513) );
  NAND2_X1 U565 ( .A1(n528), .A2(n513), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(n507), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n513), .A2(n531), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n508), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n509), .ZN(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n511) );
  NAND2_X1 U572 ( .A1(n542), .A2(n513), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n537), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U577 ( .A1(n577), .A2(n563), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n515), .A2(n526), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(n516), .Z(n523) );
  NAND2_X1 U580 ( .A1(n523), .A2(n528), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n531), .A2(n523), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(n521), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n542), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U590 ( .A1(n523), .A2(n537), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  XOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT109), .Z(n530) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n538), .A2(n528), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1336GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n533) );
  NAND2_X1 U597 ( .A1(n538), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n542), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(KEYINPUT112), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G99GAT), .B(n536), .ZN(G1338GAT) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(KEYINPUT44), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n557), .A2(n543), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n560), .A2(n552), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n544), .B(KEYINPUT114), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U612 ( .A1(n552), .A2(n563), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n549) );
  NAND2_X1 U615 ( .A1(n552), .A2(n587), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G134GAT), .B(n555), .ZN(G1343GAT) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n575), .A2(n558), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT117), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n560), .A2(n571), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT118), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U629 ( .A1(n571), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT119), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n571), .A2(n587), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT120), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n569), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n587), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n590) );
  NOR2_X1 U641 ( .A1(n577), .A2(n590), .ZN(n582) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT124), .B(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U648 ( .A(n590), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n588), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n498), .A2(n590), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

