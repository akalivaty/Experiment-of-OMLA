

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801;

  AND2_X1 U375 ( .A1(n474), .A2(n476), .ZN(n357) );
  AND2_X1 U376 ( .A1(n657), .A2(n683), .ZN(n469) );
  XNOR2_X1 U377 ( .A(n371), .B(KEYINPUT89), .ZN(n375) );
  AND2_X1 U378 ( .A1(n413), .A2(n409), .ZN(n440) );
  NAND2_X1 U379 ( .A1(n456), .A2(n459), .ZN(n371) );
  AND2_X1 U380 ( .A1(n463), .A2(n385), .ZN(n456) );
  XNOR2_X1 U381 ( .A(n360), .B(G119), .ZN(n408) );
  XNOR2_X2 U382 ( .A(n381), .B(n524), .ZN(n690) );
  NAND2_X1 U383 ( .A1(n799), .A2(n800), .ZN(n475) );
  XNOR2_X2 U384 ( .A(n382), .B(KEYINPUT40), .ZN(n800) );
  XNOR2_X2 U385 ( .A(n358), .B(n356), .ZN(n428) );
  NOR2_X2 U386 ( .A1(n685), .A2(n391), .ZN(n433) );
  BUF_X2 U387 ( .A(n656), .Z(n657) );
  INV_X1 U388 ( .A(n440), .ZN(n362) );
  XNOR2_X1 U389 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n356) );
  OR2_X1 U390 ( .A1(n380), .A2(n460), .ZN(n459) );
  INV_X2 U391 ( .A(G953), .ZN(n791) );
  XNOR2_X1 U392 ( .A(n642), .B(n641), .ZN(n649) );
  NAND2_X1 U393 ( .A1(n384), .A2(n465), .ZN(n358) );
  AND2_X1 U394 ( .A1(n396), .A2(n362), .ZN(n467) );
  XNOR2_X1 U395 ( .A(n376), .B(KEYINPUT0), .ZN(n384) );
  XNOR2_X1 U396 ( .A(n408), .B(n363), .ZN(n772) );
  INV_X1 U397 ( .A(KEYINPUT4), .ZN(n367) );
  XNOR2_X1 U398 ( .A(n648), .B(n647), .ZN(n425) );
  XNOR2_X1 U399 ( .A(n486), .B(n485), .ZN(n798) );
  XNOR2_X1 U400 ( .A(n643), .B(KEYINPUT104), .ZN(n685) );
  XNOR2_X1 U401 ( .A(n577), .B(n434), .ZN(n612) );
  AND2_X1 U402 ( .A1(n649), .A2(n467), .ZN(n643) );
  AND2_X1 U403 ( .A1(n649), .A2(n362), .ZN(n361) );
  OR2_X1 U404 ( .A1(n600), .A2(n579), .ZN(n577) );
  XNOR2_X1 U405 ( .A(n401), .B(n373), .ZN(n372) );
  NOR2_X1 U406 ( .A1(n364), .A2(n625), .ZN(n400) );
  NOR2_X1 U407 ( .A1(n528), .A2(n583), .ZN(n432) );
  XNOR2_X1 U408 ( .A(n371), .B(n365), .ZN(n364) );
  AND2_X1 U409 ( .A1(n482), .A2(n481), .ZN(n480) );
  NAND2_X1 U410 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X1 U411 ( .A(n772), .B(n570), .ZN(n402) );
  XNOR2_X1 U412 ( .A(n522), .B(n521), .ZN(n524) );
  XNOR2_X1 U413 ( .A(n359), .B(n519), .ZN(n522) );
  XNOR2_X1 U414 ( .A(n408), .B(n517), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n569), .B(n517), .ZN(n363) );
  XNOR2_X1 U416 ( .A(G119), .B(KEYINPUT23), .ZN(n532) );
  XNOR2_X1 U417 ( .A(KEYINPUT89), .B(KEYINPUT19), .ZN(n365) );
  XNOR2_X1 U418 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  INV_X1 U419 ( .A(n428), .ZN(n725) );
  XNOR2_X2 U420 ( .A(G116), .B(KEYINPUT3), .ZN(n360) );
  NAND2_X1 U421 ( .A1(n523), .A2(KEYINPUT4), .ZN(n368) );
  NAND2_X1 U422 ( .A1(n366), .A2(n367), .ZN(n369) );
  NAND2_X1 U423 ( .A1(n368), .A2(n369), .ZN(n784) );
  INV_X1 U424 ( .A(n523), .ZN(n366) );
  AND2_X2 U425 ( .A1(n471), .A2(n470), .ZN(n370) );
  AND2_X2 U426 ( .A1(n471), .A2(n470), .ZN(n702) );
  NOR2_X2 U427 ( .A1(n626), .A2(n730), .ZN(n627) );
  INV_X1 U428 ( .A(n372), .ZN(n756) );
  XOR2_X1 U429 ( .A(n628), .B(KEYINPUT33), .Z(n373) );
  XNOR2_X1 U430 ( .A(n375), .B(KEYINPUT19), .ZN(n374) );
  NOR2_X1 U431 ( .A1(n374), .A2(n625), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n531), .ZN(n538) );
  NAND2_X1 U433 ( .A1(n529), .A2(G221), .ZN(n377) );
  XNOR2_X2 U434 ( .A(n530), .B(n555), .ZN(n531) );
  XNOR2_X1 U435 ( .A(n378), .B(n379), .ZN(n598) );
  NOR2_X1 U436 ( .A1(n706), .A2(G902), .ZN(n378) );
  XOR2_X1 U437 ( .A(n561), .B(KEYINPUT67), .Z(n379) );
  XNOR2_X1 U438 ( .A(n424), .B(n402), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n424), .B(n402), .ZN(n668) );
  BUF_X1 U440 ( .A(n554), .Z(n381) );
  NAND2_X1 U441 ( .A1(n605), .A2(n612), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n403), .B(n659), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n403), .B(n659), .ZN(n665) );
  XNOR2_X1 U444 ( .A(n400), .B(KEYINPUT0), .ZN(n466) );
  NOR2_X1 U445 ( .A1(n464), .A2(n388), .ZN(n481) );
  NOR2_X1 U446 ( .A1(n667), .A2(n666), .ZN(n766) );
  NOR2_X1 U447 ( .A1(G953), .A2(G237), .ZN(n520) );
  NAND2_X1 U448 ( .A1(n660), .A2(n451), .ZN(n449) );
  NOR2_X1 U449 ( .A1(n633), .A2(n431), .ZN(n430) );
  XNOR2_X1 U450 ( .A(n475), .B(n591), .ZN(n474) );
  XNOR2_X1 U451 ( .A(n484), .B(n527), .ZN(n528) );
  NAND2_X1 U452 ( .A1(n480), .A2(n479), .ZN(n484) );
  OR2_X1 U453 ( .A1(n690), .A2(n423), .ZN(n422) );
  XOR2_X1 U454 ( .A(KEYINPUT100), .B(KEYINPUT5), .Z(n518) );
  XNOR2_X1 U455 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n444) );
  XNOR2_X1 U456 ( .A(G122), .B(G113), .ZN(n493) );
  XOR2_X1 U457 ( .A(KEYINPUT12), .B(G140), .Z(n494) );
  XNOR2_X1 U458 ( .A(n442), .B(G131), .ZN(n441) );
  NAND2_X1 U459 ( .A1(n520), .A2(G214), .ZN(n442) );
  XNOR2_X1 U460 ( .A(n455), .B(n454), .ZN(n664) );
  INV_X1 U461 ( .A(KEYINPUT48), .ZN(n454) );
  NAND2_X1 U462 ( .A1(n357), .A2(n477), .ZN(n455) );
  XNOR2_X1 U463 ( .A(n478), .B(KEYINPUT81), .ZN(n477) );
  NAND2_X1 U464 ( .A1(n461), .A2(n660), .ZN(n460) );
  INV_X1 U465 ( .A(n575), .ZN(n461) );
  INV_X1 U466 ( .A(n420), .ZN(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n506) );
  XOR2_X1 U468 ( .A(G134), .B(KEYINPUT7), .Z(n502) );
  XNOR2_X1 U469 ( .A(n578), .B(KEYINPUT39), .ZN(n434) );
  XNOR2_X1 U470 ( .A(n446), .B(n445), .ZN(n604) );
  XNOR2_X1 U471 ( .A(n499), .B(G475), .ZN(n445) );
  OR2_X1 U472 ( .A1(n677), .A2(G902), .ZN(n446) );
  AND2_X1 U473 ( .A1(n603), .A2(n604), .ZN(n605) );
  NOR2_X1 U474 ( .A1(n766), .A2(n390), .ZN(n437) );
  INV_X1 U475 ( .A(G237), .ZN(n526) );
  XOR2_X1 U476 ( .A(G140), .B(G137), .Z(n555) );
  XNOR2_X1 U477 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n565) );
  NAND2_X1 U478 ( .A1(G237), .A2(G234), .ZN(n511) );
  XNOR2_X1 U479 ( .A(n438), .B(KEYINPUT107), .ZN(n614) );
  AND2_X1 U480 ( .A1(n722), .A2(n439), .ZN(n438) );
  AND2_X1 U481 ( .A1(n440), .A2(n593), .ZN(n439) );
  XNOR2_X1 U482 ( .A(n559), .B(n387), .ZN(n521) );
  INV_X1 U483 ( .A(G104), .ZN(n552) );
  XNOR2_X1 U484 ( .A(KEYINPUT16), .B(G122), .ZN(n569) );
  XNOR2_X1 U485 ( .A(G128), .B(G110), .ZN(n535) );
  XNOR2_X1 U486 ( .A(n443), .B(n441), .ZN(n498) );
  XNOR2_X1 U487 ( .A(n491), .B(n444), .ZN(n443) );
  AND2_X2 U488 ( .A1(n664), .A2(n620), .ZN(n789) );
  BUF_X1 U489 ( .A(n582), .Z(n733) );
  NAND2_X1 U490 ( .A1(n412), .A2(n410), .ZN(n409) );
  NOR2_X1 U491 ( .A1(n411), .A2(n594), .ZN(n410) );
  BUF_X1 U492 ( .A(n626), .Z(n731) );
  XNOR2_X1 U493 ( .A(n509), .B(n508), .ZN(n686) );
  XNOR2_X1 U494 ( .A(n677), .B(KEYINPUT59), .ZN(n678) );
  XNOR2_X1 U495 ( .A(n380), .B(n670), .ZN(n671) );
  XNOR2_X1 U496 ( .A(n673), .B(KEYINPUT91), .ZN(n709) );
  INV_X1 U497 ( .A(n741), .ZN(n465) );
  INV_X1 U498 ( .A(KEYINPUT111), .ZN(n485) );
  INV_X1 U499 ( .A(n611), .ZN(n720) );
  INV_X1 U500 ( .A(G101), .ZN(n769) );
  NAND2_X1 U501 ( .A1(n436), .A2(n435), .ZN(n768) );
  NOR2_X1 U502 ( .A1(n767), .A2(n389), .ZN(n435) );
  NAND2_X1 U503 ( .A1(n765), .A2(n437), .ZN(n436) );
  NOR2_X1 U504 ( .A1(n458), .A2(n464), .ZN(n385) );
  XOR2_X1 U505 ( .A(n770), .B(KEYINPUT69), .Z(n386) );
  AND2_X1 U506 ( .A1(n520), .A2(G210), .ZN(n387) );
  AND2_X1 U507 ( .A1(n585), .A2(G902), .ZN(n388) );
  OR2_X1 U508 ( .A1(n729), .A2(G953), .ZN(n389) );
  AND2_X1 U509 ( .A1(n666), .A2(n764), .ZN(n390) );
  AND2_X1 U510 ( .A1(n427), .A2(n637), .ZN(n391) );
  AND2_X1 U511 ( .A1(n604), .A2(n601), .ZN(n392) );
  NOR2_X1 U512 ( .A1(n749), .A2(n640), .ZN(n393) );
  NOR2_X1 U513 ( .A1(n635), .A2(n634), .ZN(n394) );
  AND2_X1 U514 ( .A1(n459), .A2(n462), .ZN(n395) );
  INV_X1 U515 ( .A(G902), .ZN(n539) );
  AND2_X1 U516 ( .A1(n731), .A2(n733), .ZN(n396) );
  NOR2_X1 U517 ( .A1(n611), .A2(n610), .ZN(n397) );
  INV_X1 U518 ( .A(n746), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n398) );
  BUF_X1 U520 ( .A(n697), .Z(n399) );
  XNOR2_X2 U521 ( .A(n567), .B(KEYINPUT10), .ZN(n530) );
  XNOR2_X1 U522 ( .A(n706), .B(n705), .ZN(n707) );
  BUF_X1 U523 ( .A(n598), .Z(n634) );
  XNOR2_X1 U524 ( .A(n598), .B(KEYINPUT1), .ZN(n626) );
  NAND2_X1 U525 ( .A1(n585), .A2(G902), .ZN(n421) );
  NOR2_X1 U526 ( .A1(n585), .A2(G902), .ZN(n483) );
  NAND2_X1 U527 ( .A1(n627), .A2(n440), .ZN(n401) );
  INV_X1 U528 ( .A(KEYINPUT85), .ZN(n451) );
  XNOR2_X2 U529 ( .A(n554), .B(n386), .ZN(n424) );
  XNOR2_X2 U530 ( .A(n784), .B(n769), .ZN(n554) );
  NAND2_X1 U531 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U532 ( .A(n407), .B(n644), .ZN(n404) );
  NAND2_X1 U533 ( .A1(n406), .A2(n658), .ZN(n405) );
  NAND2_X1 U534 ( .A1(n468), .A2(n633), .ZN(n406) );
  NAND2_X1 U535 ( .A1(n433), .A2(n638), .ZN(n407) );
  NAND2_X1 U536 ( .A1(n412), .A2(n418), .ZN(n651) );
  INV_X1 U537 ( .A(n418), .ZN(n411) );
  INV_X1 U538 ( .A(n414), .ZN(n413) );
  NAND2_X1 U539 ( .A1(n417), .A2(n415), .ZN(n414) );
  INV_X1 U540 ( .A(n416), .ZN(n415) );
  NOR2_X1 U541 ( .A1(n418), .A2(KEYINPUT6), .ZN(n416) );
  NAND2_X1 U542 ( .A1(n420), .A2(n594), .ZN(n417) );
  NAND2_X1 U543 ( .A1(n690), .A2(n419), .ZN(n418) );
  NOR2_X1 U544 ( .A1(n585), .A2(G902), .ZN(n419) );
  INV_X1 U545 ( .A(n585), .ZN(n423) );
  XNOR2_X1 U546 ( .A(n424), .B(n560), .ZN(n706) );
  NAND2_X1 U547 ( .A1(n469), .A2(n425), .ZN(n468) );
  NAND2_X1 U548 ( .A1(n430), .A2(n425), .ZN(n658) );
  XNOR2_X1 U549 ( .A(n425), .B(G119), .ZN(G21) );
  INV_X1 U550 ( .A(n426), .ZN(n587) );
  XNOR2_X1 U551 ( .A(KEYINPUT28), .B(n586), .ZN(n426) );
  NAND2_X1 U552 ( .A1(n665), .A2(n451), .ZN(n450) );
  NAND2_X1 U553 ( .A1(n428), .A2(n636), .ZN(n427) );
  XNOR2_X1 U554 ( .A(n429), .B(n689), .ZN(G63) );
  NAND2_X1 U555 ( .A1(n688), .A2(n709), .ZN(n429) );
  INV_X1 U556 ( .A(n683), .ZN(n431) );
  NAND2_X1 U557 ( .A1(n551), .A2(n432), .ZN(n562) );
  INV_X1 U558 ( .A(n614), .ZN(n596) );
  NOR2_X1 U559 ( .A1(n789), .A2(KEYINPUT2), .ZN(n763) );
  NAND2_X1 U560 ( .A1(n627), .A2(n737), .ZN(n741) );
  NAND2_X1 U561 ( .A1(n447), .A2(n789), .ZN(n473) );
  NOR2_X1 U562 ( .A1(n452), .A2(n448), .ZN(n447) );
  NAND2_X1 U563 ( .A1(n450), .A2(n449), .ZN(n448) );
  NOR2_X1 U564 ( .A1(n383), .A2(n453), .ZN(n452) );
  NAND2_X1 U565 ( .A1(n571), .A2(KEYINPUT85), .ZN(n453) );
  INV_X2 U566 ( .A(G125), .ZN(n492) );
  NOR2_X1 U567 ( .A1(n562), .A2(n634), .ZN(n563) );
  XNOR2_X2 U568 ( .A(n492), .B(G146), .ZN(n567) );
  XNOR2_X2 U569 ( .A(n457), .B(G143), .ZN(n523) );
  XNOR2_X2 U570 ( .A(G128), .B(KEYINPUT64), .ZN(n457) );
  NAND2_X1 U571 ( .A1(n395), .A2(n463), .ZN(n595) );
  INV_X1 U572 ( .A(n462), .ZN(n458) );
  NAND2_X1 U573 ( .A1(n575), .A2(n571), .ZN(n462) );
  NAND2_X1 U574 ( .A1(n668), .A2(n575), .ZN(n463) );
  NAND2_X1 U575 ( .A1(n372), .A2(n466), .ZN(n630) );
  NAND2_X1 U576 ( .A1(n466), .A2(n393), .ZN(n642) );
  NAND2_X1 U577 ( .A1(n384), .A2(n394), .ZN(n636) );
  INV_X1 U578 ( .A(n766), .ZN(n470) );
  NAND2_X1 U579 ( .A1(n472), .A2(n489), .ZN(n471) );
  XNOR2_X1 U580 ( .A(n473), .B(KEYINPUT84), .ZN(n472) );
  NOR2_X1 U581 ( .A1(n727), .A2(n397), .ZN(n476) );
  NAND2_X1 U582 ( .A1(n608), .A2(n607), .ZN(n478) );
  OR2_X1 U583 ( .A1(n690), .A2(n423), .ZN(n479) );
  NAND2_X1 U584 ( .A1(n690), .A2(n483), .ZN(n482) );
  NAND2_X1 U585 ( .A1(n487), .A2(n392), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n488), .B(KEYINPUT110), .ZN(n487) );
  NOR2_X1 U587 ( .A1(n600), .A2(n595), .ZN(n488) );
  OR2_X1 U588 ( .A1(n660), .A2(n764), .ZN(n489) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(n587), .Z(n490) );
  INV_X1 U590 ( .A(KEYINPUT46), .ZN(n591) );
  XNOR2_X1 U591 ( .A(KEYINPUT71), .B(KEYINPUT87), .ZN(n578) );
  INV_X1 U592 ( .A(KEYINPUT60), .ZN(n681) );
  XNOR2_X1 U593 ( .A(G143), .B(G104), .ZN(n491) );
  INV_X1 U594 ( .A(n530), .ZN(n496) );
  XNOR2_X1 U595 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U596 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n498), .B(n497), .ZN(n677) );
  INV_X1 U598 ( .A(KEYINPUT13), .ZN(n499) );
  XNOR2_X1 U599 ( .A(G107), .B(G116), .ZN(n500) );
  XNOR2_X1 U600 ( .A(n500), .B(KEYINPUT103), .ZN(n504) );
  XNOR2_X1 U601 ( .A(G122), .B(KEYINPUT9), .ZN(n501) );
  XNOR2_X1 U602 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U603 ( .A(n504), .B(n503), .Z(n509) );
  NAND2_X1 U604 ( .A1(G234), .A2(n791), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n529) );
  NAND2_X1 U606 ( .A1(G217), .A2(n529), .ZN(n507) );
  XNOR2_X1 U607 ( .A(n523), .B(n507), .ZN(n508) );
  NAND2_X1 U608 ( .A1(n686), .A2(n539), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n510), .B(G478), .ZN(n601) );
  INV_X1 U610 ( .A(n601), .ZN(n603) );
  XNOR2_X1 U611 ( .A(n511), .B(KEYINPUT14), .ZN(n513) );
  NAND2_X1 U612 ( .A1(G952), .A2(n513), .ZN(n512) );
  XOR2_X1 U613 ( .A(KEYINPUT95), .B(n512), .Z(n762) );
  NOR2_X1 U614 ( .A1(n762), .A2(G953), .ZN(n624) );
  NAND2_X1 U615 ( .A1(G902), .A2(n513), .ZN(n621) );
  NOR2_X1 U616 ( .A1(G900), .A2(n621), .ZN(n514) );
  NAND2_X1 U617 ( .A1(G953), .A2(n514), .ZN(n515) );
  XOR2_X1 U618 ( .A(KEYINPUT106), .B(n515), .Z(n516) );
  NOR2_X1 U619 ( .A1(n624), .A2(n516), .ZN(n583) );
  XNOR2_X1 U620 ( .A(G113), .B(KEYINPUT92), .ZN(n517) );
  XNOR2_X1 U621 ( .A(n518), .B(G137), .ZN(n519) );
  XNOR2_X1 U622 ( .A(G134), .B(G131), .ZN(n787) );
  XNOR2_X1 U623 ( .A(n787), .B(G146), .ZN(n559) );
  INV_X1 U624 ( .A(KEYINPUT72), .ZN(n525) );
  XNOR2_X1 U625 ( .A(n525), .B(G472), .ZN(n585) );
  NAND2_X1 U626 ( .A1(n539), .A2(n526), .ZN(n572) );
  NAND2_X1 U627 ( .A1(n572), .A2(G214), .ZN(n746) );
  XOR2_X1 U628 ( .A(KEYINPUT109), .B(KEYINPUT30), .Z(n527) );
  INV_X1 U629 ( .A(n531), .ZN(n786) );
  XOR2_X1 U630 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n533) );
  XNOR2_X1 U631 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U632 ( .A(n534), .B(KEYINPUT24), .Z(n536) );
  XNOR2_X1 U633 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U634 ( .A(n538), .B(n537), .ZN(n697) );
  NAND2_X1 U635 ( .A1(n697), .A2(n539), .ZN(n544) );
  NAND2_X1 U636 ( .A1(n660), .A2(G234), .ZN(n540) );
  XNOR2_X1 U637 ( .A(n540), .B(KEYINPUT20), .ZN(n545) );
  NAND2_X1 U638 ( .A1(n545), .A2(G217), .ZN(n542) );
  XOR2_X1 U639 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n541) );
  XNOR2_X1 U640 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X2 U641 ( .A(n544), .B(n543), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n545), .A2(G221), .ZN(n547) );
  INV_X1 U643 ( .A(KEYINPUT21), .ZN(n546) );
  XNOR2_X1 U644 ( .A(n547), .B(n546), .ZN(n734) );
  INV_X1 U645 ( .A(KEYINPUT99), .ZN(n548) );
  XNOR2_X1 U646 ( .A(n734), .B(n548), .ZN(n639) );
  NAND2_X1 U647 ( .A1(n582), .A2(n639), .ZN(n550) );
  INV_X1 U648 ( .A(KEYINPUT65), .ZN(n549) );
  XNOR2_X2 U649 ( .A(n550), .B(n549), .ZN(n730) );
  INV_X1 U650 ( .A(n730), .ZN(n551) );
  XNOR2_X1 U651 ( .A(G110), .B(G107), .ZN(n553) );
  XNOR2_X1 U652 ( .A(n553), .B(n552), .ZN(n770) );
  XNOR2_X1 U653 ( .A(KEYINPUT96), .B(n555), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n791), .A2(G227), .ZN(n556) );
  XNOR2_X1 U655 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U656 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U657 ( .A(KEYINPUT68), .B(G469), .ZN(n561) );
  XNOR2_X1 U658 ( .A(n563), .B(KEYINPUT75), .ZN(n600) );
  XNOR2_X1 U659 ( .A(KEYINPUT38), .B(KEYINPUT74), .ZN(n576) );
  NAND2_X1 U660 ( .A1(n791), .A2(G224), .ZN(n564) );
  XNOR2_X1 U661 ( .A(n564), .B(KEYINPUT93), .ZN(n566) );
  XNOR2_X1 U662 ( .A(n566), .B(n565), .ZN(n568) );
  XNOR2_X1 U663 ( .A(n568), .B(n567), .ZN(n570) );
  INV_X1 U664 ( .A(n660), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n572), .A2(G210), .ZN(n574) );
  XNOR2_X1 U666 ( .A(KEYINPUT78), .B(KEYINPUT94), .ZN(n573) );
  XNOR2_X1 U667 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U668 ( .A(n576), .B(n595), .Z(n579) );
  INV_X1 U669 ( .A(n579), .ZN(n747) );
  NAND2_X1 U670 ( .A1(n747), .A2(n746), .ZN(n751) );
  INV_X1 U671 ( .A(n604), .ZN(n580) );
  NAND2_X1 U672 ( .A1(n580), .A2(n603), .ZN(n749) );
  NOR2_X1 U673 ( .A1(n751), .A2(n749), .ZN(n581) );
  XNOR2_X1 U674 ( .A(n581), .B(KEYINPUT41), .ZN(n745) );
  NOR2_X1 U675 ( .A1(n582), .A2(n583), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n584), .A2(n734), .ZN(n592) );
  NOR2_X1 U677 ( .A1(n592), .A2(n651), .ZN(n586) );
  INV_X1 U678 ( .A(n634), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n490), .A2(n588), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n745), .A2(n602), .ZN(n590) );
  XNOR2_X1 U681 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n589) );
  XNOR2_X1 U682 ( .A(n590), .B(n589), .ZN(n799) );
  INV_X1 U683 ( .A(n592), .ZN(n593) );
  XOR2_X1 U684 ( .A(KEYINPUT105), .B(n605), .Z(n722) );
  INV_X1 U685 ( .A(KEYINPUT6), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n596), .A2(n375), .ZN(n597) );
  XNOR2_X1 U687 ( .A(n597), .B(KEYINPUT36), .ZN(n599) );
  NOR2_X1 U688 ( .A1(n599), .A2(n731), .ZN(n727) );
  XNOR2_X1 U689 ( .A(n798), .B(KEYINPUT82), .ZN(n608) );
  OR2_X1 U690 ( .A1(n374), .A2(n602), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n724) );
  NOR2_X1 U692 ( .A1(n724), .A2(n605), .ZN(n752) );
  INV_X1 U693 ( .A(n752), .ZN(n637) );
  NAND2_X1 U694 ( .A1(n720), .A2(n637), .ZN(n606) );
  NAND2_X1 U695 ( .A1(n606), .A2(KEYINPUT47), .ZN(n607) );
  NOR2_X1 U696 ( .A1(KEYINPUT47), .A2(n752), .ZN(n609) );
  XNOR2_X1 U697 ( .A(n609), .B(KEYINPUT73), .ZN(n610) );
  NAND2_X1 U698 ( .A1(n724), .A2(n612), .ZN(n613) );
  XOR2_X1 U699 ( .A(KEYINPUT114), .B(n613), .Z(n801) );
  NOR2_X1 U700 ( .A1(n614), .A2(n464), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n615), .A2(n731), .ZN(n617) );
  XNOR2_X1 U702 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n616) );
  XNOR2_X1 U703 ( .A(n617), .B(n616), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n618), .A2(n595), .ZN(n684) );
  INV_X1 U705 ( .A(n684), .ZN(n619) );
  NOR2_X1 U706 ( .A1(n801), .A2(n619), .ZN(n620) );
  NOR2_X1 U707 ( .A1(G898), .A2(n791), .ZN(n773) );
  INV_X1 U708 ( .A(n773), .ZN(n622) );
  NOR2_X1 U709 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U711 ( .A(KEYINPUT70), .ZN(n628) );
  INV_X1 U712 ( .A(KEYINPUT34), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n631), .A2(n392), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(n398), .ZN(n656) );
  INV_X1 U716 ( .A(KEYINPUT44), .ZN(n633) );
  OR2_X2 U717 ( .A1(n656), .A2(n633), .ZN(n638) );
  INV_X1 U718 ( .A(n651), .ZN(n737) );
  OR2_X1 U719 ( .A1(n737), .A2(n730), .ZN(n635) );
  INV_X1 U720 ( .A(n636), .ZN(n713) );
  INV_X1 U721 ( .A(n639), .ZN(n640) );
  INV_X1 U722 ( .A(KEYINPUT22), .ZN(n641) );
  INV_X1 U723 ( .A(KEYINPUT88), .ZN(n644) );
  INV_X1 U724 ( .A(n731), .ZN(n653) );
  INV_X1 U725 ( .A(n733), .ZN(n650) );
  AND2_X1 U726 ( .A1(n653), .A2(n650), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n361), .A2(n645), .ZN(n648) );
  INV_X1 U728 ( .A(KEYINPUT77), .ZN(n646) );
  XNOR2_X1 U729 ( .A(n646), .B(KEYINPUT32), .ZN(n647) );
  INV_X1 U730 ( .A(n649), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  OR2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  OR2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n683) );
  INV_X1 U734 ( .A(KEYINPUT45), .ZN(n659) );
  INV_X1 U735 ( .A(KEYINPUT2), .ZN(n764) );
  OR2_X1 U736 ( .A1(n801), .A2(n764), .ZN(n661) );
  XNOR2_X1 U737 ( .A(KEYINPUT79), .B(n661), .ZN(n662) );
  AND2_X1 U738 ( .A1(n662), .A2(n684), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n667) );
  BUF_X1 U740 ( .A(n383), .Z(n666) );
  NAND2_X1 U741 ( .A1(n370), .A2(G210), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT80), .B(KEYINPUT54), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n669), .B(KEYINPUT55), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n672), .B(n671), .ZN(n674) );
  NOR2_X1 U745 ( .A1(n791), .A2(G952), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n674), .A2(n709), .ZN(n676) );
  INV_X1 U747 ( .A(KEYINPUT56), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n676), .B(n675), .ZN(G51) );
  NAND2_X1 U749 ( .A1(n702), .A2(G475), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n680), .A2(n709), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n682), .B(n681), .ZN(G60) );
  XNOR2_X1 U753 ( .A(n683), .B(G110), .ZN(G12) );
  XNOR2_X1 U754 ( .A(n684), .B(G140), .ZN(G42) );
  XNOR2_X1 U755 ( .A(n685), .B(n769), .ZN(G3) );
  INV_X1 U756 ( .A(KEYINPUT122), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n370), .A2(G478), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n657), .B(G122), .ZN(G24) );
  NAND2_X1 U760 ( .A1(n702), .A2(G472), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n690), .B(KEYINPUT62), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n693), .A2(n709), .ZN(n695) );
  XNOR2_X1 U764 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n694) );
  XNOR2_X1 U765 ( .A(n695), .B(n694), .ZN(G57) );
  NAND2_X1 U766 ( .A1(n370), .A2(G217), .ZN(n699) );
  XNOR2_X1 U767 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n399), .B(n696), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n699), .B(n698), .ZN(n701) );
  INV_X1 U770 ( .A(n709), .ZN(n700) );
  NOR2_X1 U771 ( .A1(n701), .A2(n700), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n702), .A2(G469), .ZN(n708) );
  XOR2_X1 U773 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n704) );
  XNOR2_X1 U774 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n703) );
  XNOR2_X1 U775 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U776 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(n711), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U779 ( .A1(n713), .A2(n722), .ZN(n712) );
  XNOR2_X1 U780 ( .A(n712), .B(G104), .ZN(G6) );
  XOR2_X1 U781 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n715) );
  NAND2_X1 U782 ( .A1(n713), .A2(n724), .ZN(n714) );
  XNOR2_X1 U783 ( .A(n715), .B(n714), .ZN(n717) );
  XOR2_X1 U784 ( .A(G107), .B(KEYINPUT26), .Z(n716) );
  XNOR2_X1 U785 ( .A(n717), .B(n716), .ZN(G9) );
  XOR2_X1 U786 ( .A(G128), .B(KEYINPUT29), .Z(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n724), .ZN(n718) );
  XNOR2_X1 U788 ( .A(n719), .B(n718), .ZN(G30) );
  NAND2_X1 U789 ( .A1(n720), .A2(n722), .ZN(n721) );
  XNOR2_X1 U790 ( .A(n721), .B(G146), .ZN(G48) );
  NAND2_X1 U791 ( .A1(n725), .A2(n722), .ZN(n723) );
  XNOR2_X1 U792 ( .A(n723), .B(G113), .ZN(G15) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U794 ( .A(n726), .B(G116), .ZN(G18) );
  XNOR2_X1 U795 ( .A(n727), .B(G125), .ZN(n728) );
  XNOR2_X1 U796 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U797 ( .A1(n745), .A2(n756), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U799 ( .A(n732), .B(KEYINPUT50), .ZN(n739) );
  NOR2_X1 U800 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U801 ( .A(KEYINPUT49), .B(n735), .Z(n736) );
  NOR2_X1 U802 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U803 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U804 ( .A(n740), .B(KEYINPUT116), .ZN(n742) );
  NAND2_X1 U805 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U806 ( .A(KEYINPUT51), .B(n743), .ZN(n744) );
  NOR2_X1 U807 ( .A1(n745), .A2(n744), .ZN(n759) );
  NOR2_X1 U808 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U809 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U810 ( .A(KEYINPUT117), .B(n750), .Z(n754) );
  NOR2_X1 U811 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U812 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U813 ( .A(n755), .B(KEYINPUT118), .ZN(n757) );
  NOR2_X1 U814 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U815 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U816 ( .A(n760), .B(KEYINPUT52), .ZN(n761) );
  NOR2_X1 U817 ( .A1(n762), .A2(n761), .ZN(n767) );
  XNOR2_X1 U818 ( .A(n763), .B(KEYINPUT83), .ZN(n765) );
  XOR2_X1 U819 ( .A(KEYINPUT53), .B(n768), .Z(G75) );
  XNOR2_X1 U820 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(n774) );
  NOR2_X1 U822 ( .A1(n774), .A2(n773), .ZN(n782) );
  INV_X1 U823 ( .A(n666), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(n791), .ZN(n780) );
  XOR2_X1 U825 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n777) );
  NAND2_X1 U826 ( .A1(G224), .A2(G953), .ZN(n776) );
  XNOR2_X1 U827 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U828 ( .A1(n778), .A2(G898), .ZN(n779) );
  NAND2_X1 U829 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U830 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U831 ( .A(KEYINPUT126), .B(n783), .ZN(G69) );
  BUF_X1 U832 ( .A(n784), .Z(n785) );
  XNOR2_X1 U833 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U834 ( .A(n785), .B(n788), .ZN(n793) );
  XNOR2_X1 U835 ( .A(KEYINPUT127), .B(n793), .ZN(n790) );
  XNOR2_X1 U836 ( .A(n790), .B(n789), .ZN(n792) );
  NAND2_X1 U837 ( .A1(n792), .A2(n791), .ZN(n797) );
  XNOR2_X1 U838 ( .A(G227), .B(n793), .ZN(n794) );
  NAND2_X1 U839 ( .A1(n794), .A2(G900), .ZN(n795) );
  NAND2_X1 U840 ( .A1(n795), .A2(G953), .ZN(n796) );
  NAND2_X1 U841 ( .A1(n797), .A2(n796), .ZN(G72) );
  XNOR2_X1 U842 ( .A(G143), .B(n798), .ZN(G45) );
  XNOR2_X1 U843 ( .A(G137), .B(n799), .ZN(G39) );
  XNOR2_X1 U844 ( .A(G131), .B(n800), .ZN(G33) );
  XOR2_X1 U845 ( .A(G134), .B(n801), .Z(G36) );
endmodule

