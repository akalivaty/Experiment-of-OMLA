

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769;

  XNOR2_X1 U375 ( .A(n461), .B(n501), .ZN(n419) );
  AND2_X2 U376 ( .A1(n414), .A2(n411), .ZN(n410) );
  AND2_X4 U377 ( .A1(n693), .A2(n650), .ZN(n683) );
  XNOR2_X2 U378 ( .A(n649), .B(KEYINPUT83), .ZN(n693) );
  XNOR2_X2 U379 ( .A(n488), .B(n428), .ZN(n530) );
  XNOR2_X2 U380 ( .A(n427), .B(n426), .ZN(n488) );
  NAND2_X1 U381 ( .A1(n397), .A2(n394), .ZN(n636) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n498) );
  INV_X1 U383 ( .A(n493), .ZN(n583) );
  AND2_X1 U384 ( .A1(n407), .A2(n404), .ZN(n403) );
  XNOR2_X1 U385 ( .A(n486), .B(n485), .ZN(n527) );
  XNOR2_X1 U386 ( .A(n379), .B(n378), .ZN(n537) );
  XNOR2_X1 U387 ( .A(n465), .B(KEYINPUT10), .ZN(n664) );
  XNOR2_X1 U388 ( .A(KEYINPUT71), .B(G131), .ZN(n501) );
  XNOR2_X1 U389 ( .A(KEYINPUT67), .B(G101), .ZN(n463) );
  XNOR2_X1 U390 ( .A(G146), .B(G125), .ZN(n465) );
  XNOR2_X1 U391 ( .A(G143), .B(G128), .ZN(n464) );
  NAND2_X1 U392 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U393 ( .A(n549), .B(n548), .ZN(n354) );
  BUF_X1 U394 ( .A(n677), .Z(n355) );
  XNOR2_X1 U395 ( .A(n549), .B(n548), .ZN(n559) );
  NOR2_X1 U396 ( .A1(n661), .A2(n657), .ZN(n562) );
  AND2_X1 U397 ( .A1(n535), .A2(n660), .ZN(n556) );
  OR2_X1 U398 ( .A1(n751), .A2(n736), .ZN(n524) );
  NAND2_X1 U399 ( .A1(n699), .A2(n698), .ZN(n695) );
  OR2_X1 U400 ( .A1(n696), .A2(n699), .ZN(n550) );
  INV_X1 U401 ( .A(KEYINPUT0), .ZN(n485) );
  XNOR2_X1 U402 ( .A(n557), .B(KEYINPUT97), .ZN(n566) );
  NOR2_X1 U403 ( .A1(G902), .A2(G237), .ZN(n472) );
  NAND2_X1 U404 ( .A1(n396), .A2(n567), .ZN(n395) );
  INV_X1 U405 ( .A(n474), .ZN(n396) );
  XNOR2_X1 U406 ( .A(G119), .B(G116), .ZN(n451) );
  INV_X1 U407 ( .A(n689), .ZN(n406) );
  NOR2_X1 U408 ( .A1(n397), .A2(n478), .ZN(n392) );
  XNOR2_X1 U409 ( .A(n506), .B(n505), .ZN(n675) );
  XNOR2_X1 U410 ( .A(n504), .B(n416), .ZN(n505) );
  AND2_X1 U411 ( .A1(n595), .A2(n590), .ZN(n591) );
  XNOR2_X1 U412 ( .A(n529), .B(n360), .ZN(n532) );
  NOR2_X1 U413 ( .A1(n672), .A2(G902), .ZN(n375) );
  NOR2_X1 U414 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U415 ( .A(n630), .B(KEYINPUT72), .ZN(n631) );
  XNOR2_X1 U416 ( .A(n430), .B(n429), .ZN(n510) );
  XNOR2_X1 U417 ( .A(KEYINPUT99), .B(KEYINPUT17), .ZN(n460) );
  INV_X1 U418 ( .A(KEYINPUT81), .ZN(n378) );
  NOR2_X1 U419 ( .A1(n477), .A2(KEYINPUT19), .ZN(n390) );
  NAND2_X1 U420 ( .A1(n387), .A2(n386), .ZN(n393) );
  NAND2_X1 U421 ( .A1(n477), .A2(KEYINPUT19), .ZN(n386) );
  OR2_X1 U422 ( .A1(n395), .A2(n478), .ZN(n388) );
  AND2_X1 U423 ( .A1(n399), .A2(n398), .ZN(n397) );
  NAND2_X1 U424 ( .A1(n474), .A2(n644), .ZN(n398) );
  XNOR2_X1 U425 ( .A(G113), .B(KEYINPUT75), .ZN(n450) );
  XNOR2_X1 U426 ( .A(G128), .B(G119), .ZN(n435) );
  XNOR2_X1 U427 ( .A(KEYINPUT90), .B(G110), .ZN(n431) );
  XNOR2_X1 U428 ( .A(G107), .B(G116), .ZN(n511) );
  NOR2_X1 U429 ( .A1(n406), .A2(n405), .ZN(n404) );
  NOR2_X1 U430 ( .A1(n644), .A2(n569), .ZN(n405) );
  NAND2_X1 U431 ( .A1(n402), .A2(KEYINPUT92), .ZN(n401) );
  XNOR2_X1 U432 ( .A(G110), .B(G107), .ZN(n420) );
  XNOR2_X1 U433 ( .A(n571), .B(n570), .ZN(n727) );
  AND2_X1 U434 ( .A1(n415), .A2(n545), .ZN(n411) );
  NAND2_X1 U435 ( .A1(n412), .A2(n413), .ZN(n409) );
  NOR2_X1 U436 ( .A1(n581), .A2(n489), .ZN(n605) );
  BUF_X1 U437 ( .A(n530), .Z(n696) );
  XNOR2_X1 U438 ( .A(n507), .B(G475), .ZN(n508) );
  XNOR2_X1 U439 ( .A(n400), .B(KEYINPUT42), .ZN(n769) );
  NAND2_X1 U440 ( .A1(n727), .A2(n605), .ZN(n400) );
  XNOR2_X1 U441 ( .A(n592), .B(KEYINPUT40), .ZN(n768) );
  XNOR2_X1 U442 ( .A(n553), .B(n552), .ZN(n661) );
  OR2_X1 U443 ( .A1(n540), .A2(n490), .ZN(n492) );
  XNOR2_X1 U444 ( .A(n384), .B(KEYINPUT106), .ZN(n660) );
  INV_X1 U445 ( .A(KEYINPUT96), .ZN(n533) );
  INV_X1 U446 ( .A(KEYINPUT60), .ZN(n371) );
  INV_X1 U447 ( .A(KEYINPUT56), .ZN(n367) );
  XOR2_X1 U448 ( .A(n424), .B(n423), .Z(n356) );
  XOR2_X1 U449 ( .A(n443), .B(n442), .Z(n357) );
  AND2_X1 U450 ( .A1(n551), .A2(n618), .ZN(n358) );
  AND2_X1 U451 ( .A1(n394), .A2(n390), .ZN(n359) );
  XOR2_X1 U452 ( .A(n528), .B(KEYINPUT22), .Z(n360) );
  INV_X1 U453 ( .A(KEYINPUT19), .ZN(n478) );
  XOR2_X1 U454 ( .A(n652), .B(n651), .Z(n361) );
  XNOR2_X1 U455 ( .A(n675), .B(KEYINPUT59), .ZN(n362) );
  XOR2_X1 U456 ( .A(n685), .B(n684), .Z(n363) );
  AND2_X1 U457 ( .A1(n644), .A2(n569), .ZN(n364) );
  NOR2_X1 U458 ( .A1(n665), .A2(G952), .ZN(n687) );
  INV_X1 U459 ( .A(n687), .ZN(n373) );
  NAND2_X1 U460 ( .A1(n365), .A2(KEYINPUT44), .ZN(n377) );
  NAND2_X1 U461 ( .A1(n354), .A2(n562), .ZN(n365) );
  XNOR2_X1 U462 ( .A(n366), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U463 ( .A1(n369), .A2(n373), .ZN(n366) );
  XNOR2_X1 U464 ( .A(n368), .B(n367), .ZN(G51) );
  NAND2_X1 U465 ( .A1(n370), .A2(n373), .ZN(n368) );
  XNOR2_X1 U466 ( .A(n663), .B(n662), .ZN(n369) );
  XNOR2_X1 U467 ( .A(n686), .B(n363), .ZN(n370) );
  NOR2_X1 U468 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U469 ( .A(n372), .B(n371), .ZN(G60) );
  NAND2_X1 U470 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U471 ( .A1(n532), .A2(n358), .ZN(n553) );
  XNOR2_X1 U472 ( .A(n383), .B(n465), .ZN(n376) );
  XNOR2_X1 U473 ( .A(n376), .B(n466), .ZN(n382) );
  XNOR2_X1 U474 ( .A(n676), .B(n362), .ZN(n374) );
  NAND2_X1 U475 ( .A1(n510), .A2(G221), .ZN(n434) );
  XNOR2_X2 U476 ( .A(n375), .B(n357), .ZN(n699) );
  NAND2_X1 U477 ( .A1(n532), .A2(n417), .ZN(n534) );
  NOR2_X1 U478 ( .A1(n585), .A2(n586), .ZN(n588) );
  NOR2_X1 U479 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U480 ( .A1(n377), .A2(n556), .ZN(n557) );
  NOR2_X2 U481 ( .A1(n530), .A2(n695), .ZN(n379) );
  XNOR2_X1 U482 ( .A(n380), .B(n356), .ZN(n677) );
  XNOR2_X1 U483 ( .A(n380), .B(n664), .ZN(n667) );
  XNOR2_X2 U484 ( .A(n455), .B(n437), .ZN(n380) );
  XNOR2_X1 U485 ( .A(n382), .B(n381), .ZN(n471) );
  XNOR2_X1 U486 ( .A(n461), .B(n462), .ZN(n381) );
  XNOR2_X2 U487 ( .A(n418), .B(KEYINPUT4), .ZN(n461) );
  XNOR2_X1 U488 ( .A(n460), .B(KEYINPUT18), .ZN(n383) );
  NAND2_X1 U489 ( .A1(n385), .A2(n699), .ZN(n384) );
  XNOR2_X1 U490 ( .A(n534), .B(n533), .ZN(n385) );
  OR2_X1 U491 ( .A1(n685), .A2(n395), .ZN(n394) );
  OR2_X1 U492 ( .A1(n685), .A2(n388), .ZN(n387) );
  NAND2_X1 U493 ( .A1(n391), .A2(n389), .ZN(n606) );
  NAND2_X1 U494 ( .A1(n397), .A2(n359), .ZN(n389) );
  NAND2_X1 U495 ( .A1(n685), .A2(n474), .ZN(n399) );
  NAND2_X1 U496 ( .A1(n769), .A2(n768), .ZN(n593) );
  NAND2_X1 U497 ( .A1(n403), .A2(n401), .ZN(n408) );
  INV_X1 U498 ( .A(n568), .ZN(n402) );
  NAND2_X1 U499 ( .A1(n568), .A2(n364), .ZN(n407) );
  NAND2_X1 U500 ( .A1(n408), .A2(n645), .ZN(n650) );
  NAND2_X2 U501 ( .A1(n410), .A2(n409), .ZN(n549) );
  INV_X1 U502 ( .A(n717), .ZN(n412) );
  XNOR2_X2 U503 ( .A(n539), .B(n538), .ZN(n717) );
  NOR2_X1 U504 ( .A1(n540), .A2(n541), .ZN(n413) );
  NAND2_X1 U505 ( .A1(n717), .A2(n541), .ZN(n414) );
  NAND2_X1 U506 ( .A1(n540), .A2(n541), .ZN(n415) );
  XOR2_X1 U507 ( .A(n503), .B(n502), .Z(n416) );
  AND2_X1 U508 ( .A1(n696), .A2(n618), .ZN(n417) );
  NOR2_X1 U509 ( .A1(KEYINPUT69), .A2(n714), .ZN(n609) );
  XNOR2_X1 U510 ( .A(n431), .B(KEYINPUT24), .ZN(n432) );
  BUF_X1 U511 ( .A(n717), .Z(n726) );
  XNOR2_X1 U512 ( .A(n664), .B(n432), .ZN(n433) );
  XNOR2_X1 U513 ( .A(n509), .B(n508), .ZN(n542) );
  XNOR2_X2 U514 ( .A(KEYINPUT65), .B(KEYINPUT70), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n464), .B(G134), .ZN(n516) );
  XNOR2_X2 U516 ( .A(n419), .B(n516), .ZN(n455) );
  XNOR2_X1 U517 ( .A(G140), .B(G137), .ZN(n437) );
  XNOR2_X1 U518 ( .A(n463), .B(G146), .ZN(n449) );
  XNOR2_X1 U519 ( .A(n420), .B(G104), .ZN(n468) );
  XNOR2_X1 U520 ( .A(n449), .B(n468), .ZN(n424) );
  INV_X1 U521 ( .A(KEYINPUT64), .ZN(n421) );
  XNOR2_X2 U522 ( .A(n421), .B(G953), .ZN(n665) );
  NAND2_X1 U523 ( .A1(n665), .A2(G227), .ZN(n422) );
  XNOR2_X1 U524 ( .A(n422), .B(KEYINPUT85), .ZN(n423) );
  OR2_X2 U525 ( .A1(n677), .A2(G902), .ZN(n427) );
  XNOR2_X1 U526 ( .A(KEYINPUT74), .B(G469), .ZN(n425) );
  XNOR2_X1 U527 ( .A(n425), .B(KEYINPUT73), .ZN(n426) );
  XNOR2_X1 U528 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n428) );
  NAND2_X1 U529 ( .A1(n665), .A2(G234), .ZN(n430) );
  XNOR2_X1 U530 ( .A(KEYINPUT91), .B(KEYINPUT8), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n434), .B(n433), .ZN(n440) );
  XOR2_X1 U532 ( .A(KEYINPUT23), .B(KEYINPUT101), .Z(n436) );
  XNOR2_X1 U533 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U534 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U535 ( .A(n440), .B(n439), .ZN(n672) );
  XOR2_X1 U536 ( .A(KEYINPUT25), .B(KEYINPUT84), .Z(n443) );
  XNOR2_X1 U537 ( .A(KEYINPUT15), .B(G902), .ZN(n567) );
  NAND2_X1 U538 ( .A1(n567), .A2(G234), .ZN(n441) );
  XNOR2_X1 U539 ( .A(n441), .B(KEYINPUT20), .ZN(n444) );
  NAND2_X1 U540 ( .A1(n444), .A2(G217), .ZN(n442) );
  AND2_X1 U541 ( .A1(n444), .A2(G221), .ZN(n445) );
  XNOR2_X1 U542 ( .A(n445), .B(KEYINPUT21), .ZN(n698) );
  XOR2_X1 U543 ( .A(G137), .B(KEYINPUT5), .Z(n447) );
  NAND2_X1 U544 ( .A1(n498), .A2(G210), .ZN(n446) );
  XNOR2_X1 U545 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n449), .B(n448), .ZN(n454) );
  XNOR2_X1 U547 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U548 ( .A(KEYINPUT98), .B(KEYINPUT3), .ZN(n452) );
  XNOR2_X1 U549 ( .A(n453), .B(n452), .ZN(n470) );
  XNOR2_X1 U550 ( .A(n454), .B(n470), .ZN(n456) );
  XNOR2_X1 U551 ( .A(n455), .B(n456), .ZN(n652) );
  INV_X1 U552 ( .A(G902), .ZN(n519) );
  NAND2_X1 U553 ( .A1(n652), .A2(n519), .ZN(n459) );
  INV_X1 U554 ( .A(KEYINPUT78), .ZN(n457) );
  XNOR2_X1 U555 ( .A(n457), .B(G472), .ZN(n458) );
  XNOR2_X2 U556 ( .A(n459), .B(n458), .ZN(n493) );
  AND2_X1 U557 ( .A1(n537), .A2(n583), .ZN(n704) );
  NAND2_X1 U558 ( .A1(n665), .A2(G224), .ZN(n462) );
  XNOR2_X1 U559 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U560 ( .A(G122), .B(KEYINPUT16), .ZN(n467) );
  XNOR2_X1 U561 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U562 ( .A(n470), .B(n469), .ZN(n762) );
  XNOR2_X1 U563 ( .A(n471), .B(n762), .ZN(n685) );
  INV_X1 U564 ( .A(n567), .ZN(n644) );
  XNOR2_X1 U565 ( .A(n472), .B(KEYINPUT82), .ZN(n476) );
  INV_X1 U566 ( .A(G210), .ZN(n473) );
  OR2_X1 U567 ( .A1(n476), .A2(n473), .ZN(n474) );
  INV_X1 U568 ( .A(G214), .ZN(n475) );
  OR2_X1 U569 ( .A1(n476), .A2(n475), .ZN(n708) );
  INV_X1 U570 ( .A(n708), .ZN(n477) );
  NAND2_X1 U571 ( .A1(G237), .A2(G234), .ZN(n479) );
  XNOR2_X1 U572 ( .A(n479), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U573 ( .A1(G952), .A2(n481), .ZN(n480) );
  XNOR2_X1 U574 ( .A(KEYINPUT100), .B(n480), .ZN(n723) );
  NOR2_X1 U575 ( .A1(n723), .A2(G953), .ZN(n575) );
  AND2_X1 U576 ( .A1(G902), .A2(n481), .ZN(n573) );
  INV_X1 U577 ( .A(G898), .ZN(n482) );
  AND2_X1 U578 ( .A1(n482), .A2(G953), .ZN(n763) );
  AND2_X1 U579 ( .A1(n573), .A2(n763), .ZN(n483) );
  OR2_X1 U580 ( .A1(n575), .A2(n483), .ZN(n484) );
  NAND2_X1 U581 ( .A1(n606), .A2(n484), .ZN(n486) );
  NAND2_X1 U582 ( .A1(n704), .A2(n527), .ZN(n487) );
  XNOR2_X1 U583 ( .A(n487), .B(KEYINPUT31), .ZN(n751) );
  INV_X1 U584 ( .A(n527), .ZN(n540) );
  BUF_X1 U585 ( .A(n488), .Z(n489) );
  OR2_X1 U586 ( .A1(n489), .A2(n695), .ZN(n490) );
  INV_X1 U587 ( .A(KEYINPUT102), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n492), .B(n491), .ZN(n494) );
  AND2_X1 U589 ( .A1(n494), .A2(n493), .ZN(n736) );
  XOR2_X1 U590 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n496) );
  XNOR2_X1 U591 ( .A(G122), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U592 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U593 ( .A(n664), .B(n497), .Z(n500) );
  NAND2_X1 U594 ( .A1(n498), .A2(G214), .ZN(n499) );
  XNOR2_X1 U595 ( .A(n500), .B(n499), .ZN(n506) );
  XOR2_X1 U596 ( .A(KEYINPUT11), .B(n501), .Z(n504) );
  XOR2_X1 U597 ( .A(G140), .B(G113), .Z(n503) );
  XNOR2_X1 U598 ( .A(G143), .B(G104), .ZN(n502) );
  NOR2_X1 U599 ( .A1(G902), .A2(n675), .ZN(n509) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(KEYINPUT105), .ZN(n507) );
  AND2_X1 U601 ( .A1(n510), .A2(G217), .ZN(n514) );
  XNOR2_X1 U602 ( .A(n511), .B(KEYINPUT7), .ZN(n512) );
  XOR2_X1 U603 ( .A(n512), .B(KEYINPUT9), .Z(n513) );
  XNOR2_X1 U604 ( .A(n514), .B(n513), .ZN(n518) );
  INV_X1 U605 ( .A(G122), .ZN(n515) );
  XNOR2_X1 U606 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U607 ( .A(n518), .B(n517), .ZN(n662) );
  NAND2_X1 U608 ( .A1(n662), .A2(n519), .ZN(n521) );
  INV_X1 U609 ( .A(G478), .ZN(n520) );
  XNOR2_X1 U610 ( .A(n521), .B(n520), .ZN(n525) );
  INV_X1 U611 ( .A(n525), .ZN(n543) );
  AND2_X1 U612 ( .A1(n542), .A2(n543), .ZN(n750) );
  INV_X1 U613 ( .A(n750), .ZN(n522) );
  OR2_X1 U614 ( .A1(n542), .A2(n543), .ZN(n582) );
  AND2_X1 U615 ( .A1(n522), .A2(n582), .ZN(n714) );
  INV_X1 U616 ( .A(n714), .ZN(n523) );
  NAND2_X1 U617 ( .A1(n524), .A2(n523), .ZN(n535) );
  NAND2_X1 U618 ( .A1(n542), .A2(n525), .ZN(n711) );
  INV_X1 U619 ( .A(n698), .ZN(n576) );
  NOR2_X1 U620 ( .A1(n711), .A2(n576), .ZN(n526) );
  NAND2_X1 U621 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U622 ( .A(KEYINPUT79), .ZN(n528) );
  INV_X1 U623 ( .A(KEYINPUT6), .ZN(n531) );
  XNOR2_X1 U624 ( .A(n493), .B(n531), .ZN(n618) );
  INV_X1 U625 ( .A(n618), .ZN(n536) );
  INV_X1 U626 ( .A(KEYINPUT33), .ZN(n538) );
  XOR2_X1 U627 ( .A(KEYINPUT77), .B(KEYINPUT34), .Z(n541) );
  INV_X1 U628 ( .A(n542), .ZN(n544) );
  NAND2_X1 U629 ( .A1(n544), .A2(n543), .ZN(n596) );
  XNOR2_X1 U630 ( .A(n596), .B(KEYINPUT87), .ZN(n545) );
  XNOR2_X1 U631 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n547) );
  INV_X1 U632 ( .A(KEYINPUT86), .ZN(n546) );
  XNOR2_X1 U633 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U634 ( .A(n550), .B(KEYINPUT107), .ZN(n551) );
  INV_X1 U635 ( .A(KEYINPUT32), .ZN(n552) );
  INV_X1 U636 ( .A(n699), .ZN(n577) );
  AND2_X1 U637 ( .A1(n577), .A2(n493), .ZN(n554) );
  AND2_X1 U638 ( .A1(n696), .A2(n554), .ZN(n555) );
  AND2_X1 U639 ( .A1(n532), .A2(n555), .ZN(n657) );
  INV_X1 U640 ( .A(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U641 ( .A1(n559), .A2(n558), .ZN(n561) );
  INV_X1 U642 ( .A(KEYINPUT68), .ZN(n560) );
  XNOR2_X1 U643 ( .A(n561), .B(n560), .ZN(n563) );
  NAND2_X1 U644 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U645 ( .A(n564), .B(KEYINPUT76), .ZN(n565) );
  NAND2_X1 U646 ( .A1(n566), .A2(n565), .ZN(n647) );
  INV_X1 U647 ( .A(KEYINPUT45), .ZN(n646) );
  XNOR2_X1 U648 ( .A(n647), .B(KEYINPUT45), .ZN(n568) );
  INV_X1 U649 ( .A(KEYINPUT92), .ZN(n569) );
  XOR2_X1 U650 ( .A(KEYINPUT46), .B(KEYINPUT95), .Z(n594) );
  XOR2_X1 U651 ( .A(KEYINPUT38), .B(n636), .Z(n589) );
  INV_X1 U652 ( .A(n589), .ZN(n709) );
  NAND2_X1 U653 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U654 ( .A1(n711), .A2(n713), .ZN(n571) );
  XNOR2_X1 U655 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n570) );
  XOR2_X1 U656 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n580) );
  NOR2_X1 U657 ( .A1(n665), .A2(G900), .ZN(n572) );
  AND2_X1 U658 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U659 ( .A1(n575), .A2(n574), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n576), .A2(n586), .ZN(n578) );
  NAND2_X1 U661 ( .A1(n578), .A2(n577), .ZN(n617) );
  NOR2_X1 U662 ( .A1(n493), .A2(n617), .ZN(n579) );
  XNOR2_X1 U663 ( .A(n580), .B(n579), .ZN(n581) );
  INV_X1 U664 ( .A(n582), .ZN(n748) );
  NAND2_X1 U665 ( .A1(n583), .A2(n708), .ZN(n584) );
  XNOR2_X1 U666 ( .A(n584), .B(KEYINPUT30), .ZN(n585) );
  INV_X1 U667 ( .A(n695), .ZN(n587) );
  AND2_X1 U668 ( .A1(n588), .A2(n587), .ZN(n595) );
  INV_X1 U669 ( .A(n489), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n589), .A2(n489), .ZN(n590) );
  XOR2_X1 U671 ( .A(n591), .B(KEYINPUT39), .Z(n640) );
  NAND2_X1 U672 ( .A1(n748), .A2(n640), .ZN(n592) );
  XNOR2_X1 U673 ( .A(n594), .B(n593), .ZN(n629) );
  INV_X1 U674 ( .A(KEYINPUT88), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n714), .A2(KEYINPUT47), .ZN(n600) );
  INV_X1 U676 ( .A(n636), .ZN(n623) );
  NAND2_X1 U677 ( .A1(n595), .A2(n623), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n656) );
  NAND2_X1 U680 ( .A1(n600), .A2(n656), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n604), .A2(n601), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n656), .A2(KEYINPUT88), .ZN(n602) );
  AND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n615) );
  OR2_X1 U684 ( .A1(n609), .A2(n604), .ZN(n607) );
  AND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n744) );
  NAND2_X1 U686 ( .A1(n607), .A2(n744), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n608), .A2(KEYINPUT47), .ZN(n613) );
  INV_X1 U688 ( .A(n609), .ZN(n610) );
  NOR2_X1 U689 ( .A1(KEYINPUT47), .A2(n610), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n744), .A2(n611), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT80), .ZN(n627) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT108), .B(n619), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n620), .A2(n748), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT109), .ZN(n622) );
  AND2_X1 U697 ( .A1(n622), .A2(n708), .ZN(n633) );
  NAND2_X1 U698 ( .A1(n633), .A2(n623), .ZN(n624) );
  XOR2_X1 U699 ( .A(KEYINPUT36), .B(n624), .Z(n626) );
  INV_X1 U700 ( .A(n696), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n659) );
  NAND2_X1 U702 ( .A1(n627), .A2(n659), .ZN(n628) );
  INV_X1 U703 ( .A(KEYINPUT48), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n632), .B(n631), .ZN(n643) );
  NAND2_X1 U705 ( .A1(n633), .A2(n696), .ZN(n635) );
  XNOR2_X1 U706 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n639) );
  INV_X1 U709 ( .A(KEYINPUT111), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n767) );
  AND2_X1 U711 ( .A1(n640), .A2(n750), .ZN(n753) );
  INV_X1 U712 ( .A(n753), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n767), .A2(n641), .ZN(n642) );
  NOR2_X4 U714 ( .A1(n643), .A2(n642), .ZN(n689) );
  NAND2_X1 U715 ( .A1(n644), .A2(KEYINPUT2), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n688) );
  NAND2_X1 U717 ( .A1(n689), .A2(KEYINPUT2), .ZN(n648) );
  NOR2_X2 U718 ( .A1(n688), .A2(n648), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n683), .A2(G472), .ZN(n653) );
  XOR2_X1 U720 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n651) );
  XNOR2_X1 U721 ( .A(n653), .B(n361), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n654), .A2(n373), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U724 ( .A(n656), .B(G143), .ZN(G45) );
  XOR2_X1 U725 ( .A(G110), .B(n657), .Z(G12) );
  XOR2_X1 U726 ( .A(G125), .B(KEYINPUT37), .Z(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(G27) );
  XNOR2_X1 U728 ( .A(n660), .B(G101), .ZN(G3) );
  XNOR2_X1 U729 ( .A(n354), .B(G122), .ZN(G24) );
  XOR2_X1 U730 ( .A(G119), .B(n661), .Z(G21) );
  NAND2_X1 U731 ( .A1(n683), .A2(G478), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n689), .B(n667), .ZN(n666) );
  NAND2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n671) );
  INV_X1 U734 ( .A(G953), .ZN(n755) );
  XOR2_X1 U735 ( .A(G227), .B(n667), .Z(n668) );
  NAND2_X1 U736 ( .A1(n668), .A2(G900), .ZN(n669) );
  NAND2_X1 U737 ( .A1(G953), .A2(n669), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(G72) );
  NAND2_X1 U739 ( .A1(n683), .A2(G217), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n674), .A2(n687), .ZN(G66) );
  NAND2_X1 U742 ( .A1(n683), .A2(G475), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n683), .A2(G469), .ZN(n681) );
  XOR2_X1 U744 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT58), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n355), .B(n679), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n682), .A2(n687), .ZN(G54) );
  NAND2_X1 U749 ( .A1(n683), .A2(G210), .ZN(n686) );
  XOR2_X1 U750 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n684) );
  INV_X1 U751 ( .A(n688), .ZN(n756) );
  NAND2_X1 U752 ( .A1(n756), .A2(n689), .ZN(n691) );
  XNOR2_X1 U753 ( .A(KEYINPUT2), .B(KEYINPUT89), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n694), .B(KEYINPUT93), .ZN(n731) );
  NAND2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U758 ( .A(KEYINPUT50), .B(n697), .Z(n703) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U760 ( .A(n700), .B(KEYINPUT49), .ZN(n701) );
  NAND2_X1 U761 ( .A1(n493), .A2(n701), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n706), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n707), .A2(n727), .ZN(n721) );
  NOR2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U768 ( .A(KEYINPUT121), .B(n712), .Z(n716) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n718), .A2(n726), .ZN(n719) );
  XOR2_X1 U772 ( .A(KEYINPUT122), .B(n719), .Z(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U774 ( .A(KEYINPUT52), .B(n722), .Z(n724) );
  NOR2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n725), .A2(G953), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n727), .A2(n412), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n733) );
  XOR2_X1 U780 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n732) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(G75) );
  XOR2_X1 U782 ( .A(G104), .B(KEYINPUT115), .Z(n735) );
  NAND2_X1 U783 ( .A1(n736), .A2(n748), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(G6) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n738) );
  NAND2_X1 U786 ( .A1(n736), .A2(n750), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U788 ( .A(G107), .B(n739), .ZN(G9) );
  XOR2_X1 U789 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n741) );
  NAND2_X1 U790 ( .A1(n744), .A2(n750), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(n743) );
  XOR2_X1 U792 ( .A(G128), .B(KEYINPUT116), .Z(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G30) );
  XOR2_X1 U794 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n746) );
  NAND2_X1 U795 ( .A1(n744), .A2(n748), .ZN(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U797 ( .A(G146), .B(n747), .ZN(G48) );
  NAND2_X1 U798 ( .A1(n751), .A2(n748), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n749), .B(G113), .ZN(G15) );
  NAND2_X1 U800 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(G116), .ZN(G18) );
  XOR2_X1 U802 ( .A(G134), .B(n753), .Z(n754) );
  XNOR2_X1 U803 ( .A(KEYINPUT120), .B(n754), .ZN(G36) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n761) );
  NAND2_X1 U805 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U806 ( .A(n757), .B(KEYINPUT126), .ZN(n758) );
  XNOR2_X1 U807 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n766) );
  XOR2_X1 U810 ( .A(G101), .B(n762), .Z(n764) );
  NOR2_X1 U811 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n766), .B(n765), .ZN(G69) );
  XNOR2_X1 U813 ( .A(G140), .B(n767), .ZN(G42) );
  XNOR2_X1 U814 ( .A(G131), .B(n768), .ZN(G33) );
  XNOR2_X1 U815 ( .A(G137), .B(n769), .ZN(G39) );
endmodule

