//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT73), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n189), .B(new_n194), .C1(new_n190), .C2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G110), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n193), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT24), .B(G110), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT74), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(G125), .A3(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(KEYINPUT16), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n204), .B2(G140), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n208), .B2(new_n211), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n197), .B(new_n202), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G110), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n192), .A2(new_n215), .A3(new_n193), .A4(new_n195), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n200), .A2(new_n201), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n211), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  XNOR2_X1  g034(.A(G125), .B(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n209), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n214), .A2(new_n223), .A3(KEYINPUT76), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT75), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G137), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n226), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n214), .A2(new_n232), .A3(KEYINPUT76), .A4(new_n223), .ZN(new_n235));
  AOI21_X1  g049(.A(G902), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n187), .B(new_n188), .C1(new_n236), .C2(KEYINPUT77), .ZN(new_n237));
  INV_X1    g051(.A(G217), .ZN(new_n238));
  INV_X1    g052(.A(G902), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n238), .B1(G234), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n235), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n239), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT78), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT25), .B1(new_n236), .B2(new_n187), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n237), .B(new_n240), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n187), .B1(new_n236), .B2(KEYINPUT77), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(KEYINPUT25), .C1(new_n187), .C2(new_n236), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(KEYINPUT79), .A3(new_n237), .A4(new_n240), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n241), .B(KEYINPUT80), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n240), .A2(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT32), .ZN(new_n257));
  NOR2_X1   g071(.A1(G472), .A2(G902), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT31), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n209), .B2(G143), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(G128), .B1(new_n263), .B2(new_n268), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n209), .A2(G143), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G137), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n279), .A2(G134), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G137), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n277), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G131), .B1(new_n282), .B2(new_n284), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n287), .A2(KEYINPUT67), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT67), .B1(new_n287), .B2(new_n288), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT68), .B(new_n273), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n286), .B1(new_n281), .B2(new_n285), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n287), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n267), .A2(KEYINPUT0), .A3(G128), .ZN(new_n296));
  NAND2_X1  g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  OR2_X1    g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n297), .B(new_n298), .C1(new_n263), .C2(new_n271), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(new_n295), .A3(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n296), .B(new_n299), .C1(new_n303), .C2(new_n292), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n291), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n287), .A2(new_n288), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n287), .A2(KEYINPUT67), .A3(new_n288), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT68), .B1(new_n311), .B2(new_n273), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n261), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n190), .A2(G116), .ZN(new_n314));
  INV_X1    g128(.A(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT2), .B(G113), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n318), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n273), .A2(new_n288), .A3(new_n287), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n304), .A2(new_n323), .A3(KEYINPUT30), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n304), .A2(new_n323), .A3(new_n326), .A4(KEYINPUT30), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n322), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n313), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n304), .A2(new_n323), .A3(new_n322), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT26), .B(G101), .Z(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n228), .A3(G210), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n260), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g153(.A(KEYINPUT31), .B(new_n337), .C1(new_n313), .C2(new_n328), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n336), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n321), .B1(new_n306), .B2(new_n312), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(new_n330), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n330), .A2(new_n343), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n330), .A2(KEYINPUT71), .A3(new_n343), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n342), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(new_n257), .B(new_n259), .C1(new_n341), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n329), .A2(new_n338), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT31), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n329), .A2(new_n260), .A3(new_n338), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT32), .B1(new_n356), .B2(new_n258), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n336), .B1(new_n345), .B2(new_n350), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n329), .A2(new_n330), .A3(new_n342), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(KEYINPUT72), .A3(new_n349), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n304), .A2(new_n323), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n322), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(new_n364), .C1(new_n343), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n336), .A2(KEYINPUT29), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n239), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G472), .B1(new_n361), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n256), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G475), .A2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G113), .B(G122), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n206), .A2(G125), .A3(G140), .ZN(new_n378));
  AOI21_X1  g192(.A(G140), .B1(new_n206), .B2(G125), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT89), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n205), .A2(new_n381), .A3(new_n207), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(KEYINPUT19), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(KEYINPUT91), .A3(KEYINPUT19), .A4(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT19), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n221), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n385), .A2(new_n209), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n389), .A2(new_n390), .A3(new_n220), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n389), .B2(new_n220), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n332), .A2(new_n228), .A3(G214), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n262), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G131), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(KEYINPUT90), .A3(G131), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n394), .A2(G131), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n391), .A2(new_n392), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n394), .B(new_n402), .Z(new_n403));
  NAND3_X1  g217(.A1(new_n380), .A2(G146), .A3(new_n382), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n404), .A2(new_n222), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n377), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n212), .A2(new_n213), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n397), .A2(new_n399), .A3(new_n409), .A4(new_n398), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n397), .A2(new_n398), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n408), .B(new_n410), .C1(new_n411), .C2(new_n409), .ZN(new_n412));
  INV_X1    g226(.A(new_n406), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n376), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n373), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT93), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n389), .A2(new_n220), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT92), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n389), .A2(new_n390), .A3(new_n220), .ZN(new_n420));
  INV_X1    g234(.A(new_n400), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n376), .B1(new_n422), .B2(new_n413), .ZN(new_n423));
  INV_X1    g237(.A(new_n414), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n372), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT20), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n415), .A2(new_n416), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n417), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n376), .B1(new_n412), .B2(new_n413), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n239), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G475), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n433), .A2(KEYINPUT14), .A3(G116), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n433), .B2(G116), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n434), .B(new_n435), .C1(new_n315), .C2(G122), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G107), .ZN(new_n437));
  XOR2_X1   g251(.A(G116), .B(G122), .Z(new_n438));
  OR2_X1    g252(.A1(KEYINPUT81), .A2(G107), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT81), .A2(G107), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT95), .B1(new_n198), .B2(G143), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n262), .A3(G128), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n442), .A2(new_n444), .B1(new_n198), .B2(G143), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n445), .A2(new_n283), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n283), .ZN(new_n447));
  OAI221_X1 g261(.A(new_n437), .B1(new_n438), .B2(new_n441), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n438), .B(new_n441), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n450), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n442), .A2(new_n444), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n453), .A2(new_n454), .B1(new_n198), .B2(G143), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n283), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n448), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT9), .B(G234), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n459), .A2(new_n238), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n448), .B(new_n460), .C1(new_n452), .C2(new_n457), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n239), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(G478), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  AOI211_X1 g282(.A(KEYINPUT15), .B(new_n468), .C1(new_n464), .C2(new_n239), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT97), .ZN(new_n471));
  NAND2_X1  g285(.A1(G234), .A2(G237), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n472), .A2(G902), .A3(G953), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n472), .A2(G952), .A3(new_n228), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n467), .A2(new_n469), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n429), .A2(new_n432), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n209), .A2(G143), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT64), .B1(new_n262), .B2(G146), .ZN(new_n484));
  OAI211_X1 g298(.A(G128), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n198), .B1(new_n482), .B2(KEYINPUT1), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n485), .A2(KEYINPUT1), .B1(new_n486), .B2(new_n267), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT3), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n439), .A2(new_n488), .A3(G104), .A4(new_n440), .ZN(new_n489));
  INV_X1    g303(.A(G101), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n375), .A2(G107), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(KEYINPUT81), .A2(G107), .ZN(new_n494));
  NOR2_X1   g308(.A1(KEYINPUT81), .A2(G107), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n375), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n375), .A2(G107), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT10), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n488), .A2(G104), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n503), .A2(new_n494), .A3(new_n495), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n491), .A2(new_n492), .ZN(new_n505));
  OAI21_X1  g319(.A(G101), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(G101), .C1(new_n504), .C2(new_n505), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n301), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n504), .A2(new_n505), .A3(G101), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n498), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT10), .A3(new_n273), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n303), .A2(new_n292), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n502), .A2(new_n510), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G110), .B(G140), .ZN(new_n516));
  INV_X1    g330(.A(G227), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G953), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n516), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n272), .B(new_n269), .C1(new_n511), .C2(new_n498), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n500), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT84), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n500), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n294), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT12), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n530));
  NOR2_X1   g344(.A1(new_n514), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n531), .A3(KEYINPUT83), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n521), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n502), .A2(new_n510), .A3(new_n513), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n294), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n520), .B1(new_n539), .B2(new_n515), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n481), .B(new_n239), .C1(new_n537), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT85), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n538), .A2(new_n294), .ZN(new_n543));
  INV_X1    g357(.A(new_n515), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n519), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n527), .A2(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n546), .B2(new_n521), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n481), .A4(new_n239), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n500), .A2(new_n522), .A3(new_n525), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n525), .B1(new_n500), .B2(new_n522), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n550), .A2(new_n551), .A3(new_n514), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT83), .B1(new_n523), .B2(new_n531), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n523), .A2(new_n531), .A3(KEYINPUT83), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n552), .A2(KEYINPUT12), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n520), .B1(new_n555), .B2(new_n515), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n543), .A2(new_n521), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n239), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n542), .A2(new_n549), .B1(new_n558), .B2(G469), .ZN(new_n559));
  OAI21_X1  g373(.A(G221), .B1(new_n459), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G122), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g377(.A1(new_n499), .A2(new_n493), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n317), .A2(new_n318), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n314), .A2(new_n316), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT5), .ZN(new_n567));
  OAI21_X1  g381(.A(G113), .B1(new_n314), .B2(KEYINPUT5), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n563), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n572));
  AOI22_X1  g386(.A1(KEYINPUT5), .A2(new_n566), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(KEYINPUT88), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n565), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n571), .B1(new_n564), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n507), .A2(new_n321), .A3(new_n509), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n512), .A2(new_n570), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n562), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n300), .A2(G125), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n581), .A2(KEYINPUT87), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n269), .A2(new_n272), .A3(new_n204), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(KEYINPUT87), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G224), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(G953), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(KEYINPUT7), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n582), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n582), .B2(new_n584), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n580), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT86), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT6), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n506), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n321), .A2(new_n509), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n567), .A2(new_n569), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n319), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n595), .A2(new_n596), .B1(new_n564), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n562), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n579), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n603), .B2(new_n594), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n581), .A2(KEYINPUT87), .A3(new_n583), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n581), .A2(KEYINPUT87), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n586), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n582), .A2(new_n584), .A3(new_n587), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n591), .B(new_n239), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G210), .B1(G237), .B2(G902), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n594), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n602), .B2(new_n579), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n608), .B(new_n607), .C1(new_n615), .C2(new_n601), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n616), .A2(new_n239), .A3(new_n611), .A4(new_n591), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G214), .B1(G237), .B2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n559), .A2(new_n561), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n371), .A2(new_n480), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  NOR2_X1   g437(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g438(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n462), .B(new_n463), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n468), .A2(G902), .ZN(new_n628));
  INV_X1    g442(.A(new_n464), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n465), .A2(new_n468), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n429), .B2(new_n432), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n559), .A2(new_n561), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n356), .A2(new_n239), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G472), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n356), .A2(new_n258), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n256), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n620), .A2(new_n478), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n636), .A2(new_n637), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NOR2_X1   g460(.A1(new_n467), .A2(new_n469), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n432), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT20), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n426), .B1(new_n425), .B2(KEYINPUT20), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n417), .A2(KEYINPUT100), .A3(new_n427), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n428), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n653), .A2(new_n654), .A3(new_n657), .A4(new_n428), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n649), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n477), .B(KEYINPUT102), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n620), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n637), .A2(new_n659), .A3(new_n642), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NOR2_X1   g479(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n224), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n253), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n248), .A2(new_n251), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n641), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n480), .A3(new_n621), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT103), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n671), .B(new_n673), .ZN(G12));
  XOR2_X1   g488(.A(new_n475), .B(KEYINPUT104), .Z(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n473), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n669), .B1(new_n358), .B2(new_n370), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n659), .A2(new_n621), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  INV_X1    g496(.A(new_n637), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n678), .B(KEYINPUT39), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n683), .A2(KEYINPUT105), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n637), .B2(new_n684), .ZN(new_n688));
  OR3_X1    g502(.A1(new_n686), .A2(KEYINPUT40), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT40), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n429), .A2(new_n432), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n618), .B(KEYINPUT38), .Z(new_n692));
  NAND3_X1  g506(.A1(new_n248), .A2(new_n251), .A3(new_n668), .ZN(new_n693));
  INV_X1    g507(.A(new_n619), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n640), .A2(new_n257), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n259), .B1(new_n341), .B2(new_n351), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT32), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n342), .B1(new_n329), .B2(new_n330), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n366), .B2(new_n342), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n696), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n691), .A2(new_n695), .A3(new_n648), .A4(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n689), .A2(new_n690), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT106), .B(G143), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G45));
  AOI211_X1 g521(.A(new_n678), .B(new_n633), .C1(new_n429), .C2(new_n432), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n696), .A2(new_n698), .A3(new_n370), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n621), .A4(new_n693), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n712));
  INV_X1    g526(.A(new_n521), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n555), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n545), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n481), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n540), .B1(new_n555), .B2(new_n713), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT107), .B1(new_n718), .B2(G902), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n717), .A2(new_n719), .B1(new_n542), .B2(new_n549), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n712), .B1(new_n720), .B2(new_n560), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n542), .A2(new_n549), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n547), .A2(new_n716), .A3(new_n239), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(G469), .A3(new_n723), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n712), .A2(new_n722), .A3(new_n724), .A4(new_n560), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n636), .A2(new_n371), .A3(new_n643), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND4_X1  g543(.A1(new_n659), .A2(new_n371), .A3(new_n662), .A4(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  AOI21_X1  g545(.A(new_n694), .B1(new_n613), .B2(new_n617), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n560), .A2(new_n722), .A3(new_n724), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n680), .A2(KEYINPUT109), .A3(new_n480), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n709), .A2(new_n733), .A3(new_n480), .A4(new_n693), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  AOI211_X1 g553(.A(new_n647), .B(new_n620), .C1(new_n429), .C2(new_n432), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n367), .A2(new_n342), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n341), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n258), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n639), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n256), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n726), .A2(new_n660), .A3(new_n740), .A4(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT110), .B(G122), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G24));
  INV_X1    g562(.A(new_n744), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n708), .A3(new_n693), .A4(new_n733), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  OAI21_X1  g565(.A(KEYINPUT112), .B1(new_n697), .B2(KEYINPUT32), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n640), .A2(new_n753), .A3(new_n257), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(new_n754), .A3(new_n698), .A4(new_n370), .ZN(new_n755));
  INV_X1    g569(.A(new_n256), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n613), .A2(new_n619), .A3(new_n617), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n613), .A2(new_n617), .A3(KEYINPUT111), .A4(new_n619), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n763), .A2(new_n559), .A3(new_n764), .A4(new_n561), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n757), .A2(new_n758), .A3(new_n708), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n756), .A3(new_n708), .A4(new_n755), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT113), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n683), .A2(new_n763), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n371), .A3(new_n708), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n766), .A2(new_n768), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n286), .ZN(G33));
  NAND2_X1  g586(.A1(new_n656), .A2(new_n658), .ZN(new_n773));
  INV_X1    g587(.A(new_n649), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n679), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n371), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n283), .ZN(G36));
  OAI21_X1  g592(.A(new_n519), .B1(new_n546), .B2(new_n544), .ZN(new_n779));
  INV_X1    g593(.A(new_n557), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(KEYINPUT45), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT45), .B1(new_n779), .B2(new_n780), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n481), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(G469), .A2(G902), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n788), .A2(new_n789), .B1(new_n549), .B2(new_n542), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  INV_X1    g605(.A(new_n763), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n560), .A3(new_n684), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n641), .A2(new_n693), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT115), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n691), .A2(KEYINPUT43), .A3(new_n633), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT43), .B1(new_n691), .B2(new_n633), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n795), .A2(new_n800), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NAND2_X1  g618(.A1(new_n791), .A2(new_n560), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n791), .A2(KEYINPUT47), .A3(new_n560), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n709), .A2(new_n756), .A3(new_n763), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n708), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  XOR2_X1   g627(.A(new_n720), .B(KEYINPUT49), .Z(new_n814));
  NAND3_X1  g628(.A1(new_n429), .A2(new_n432), .A3(new_n632), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n692), .A2(new_n756), .A3(new_n560), .A4(new_n619), .ZN(new_n816));
  OR4_X1    g630(.A1(new_n703), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n727), .A2(new_n738), .A3(new_n730), .A4(new_n746), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n770), .A2(new_n764), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n767), .A2(KEYINPUT113), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n767), .A2(KEYINPUT113), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n777), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n647), .A2(new_n432), .A3(new_n679), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n769), .A2(new_n773), .A3(new_n680), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n634), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n691), .B2(new_n647), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n637), .A3(new_n642), .A4(new_n662), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n480), .B(new_n621), .C1(new_n371), .C2(new_n670), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n744), .A2(new_n669), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n769), .A2(new_n708), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n825), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n818), .A2(new_n822), .A3(new_n823), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n680), .A2(new_n621), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n775), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n678), .B(KEYINPUT116), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n559), .A2(new_n561), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n740), .A2(new_n669), .A3(new_n703), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n750), .A3(new_n710), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT52), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n839), .A2(new_n750), .A3(new_n710), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n681), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n834), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT117), .A3(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n847), .A2(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(KEYINPUT117), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n849), .B(new_n850), .C1(new_n834), .C2(new_n845), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT53), .B1(new_n834), .B2(new_n845), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n771), .A2(new_n832), .A3(new_n777), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n836), .A2(KEYINPUT52), .A3(new_n840), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n843), .B1(new_n842), .B2(new_n681), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n857), .A3(new_n847), .A4(new_n818), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT54), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n675), .ZN(new_n861));
  INV_X1    g675(.A(new_n720), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n561), .A3(new_n763), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n861), .A2(new_n863), .A3(new_n797), .A4(new_n796), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n757), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n703), .A2(new_n256), .A3(new_n476), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n636), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(G952), .A3(new_n228), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n796), .A2(new_n745), .A3(new_n861), .A4(new_n797), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n869), .B1(new_n733), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n692), .A2(new_n560), .A3(new_n694), .A4(new_n720), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT50), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n691), .A2(new_n632), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n867), .A2(new_n863), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n880), .A2(new_n881), .B1(new_n864), .B2(new_n830), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n862), .A2(new_n560), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n807), .A2(new_n808), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n871), .A2(new_n792), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n876), .B(new_n882), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT51), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n792), .B(new_n871), .C1(new_n809), .C2(new_n883), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n876), .A4(new_n882), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n873), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n852), .A2(new_n860), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n852), .A2(new_n860), .A3(new_n892), .A4(KEYINPUT119), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT120), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n817), .B1(new_n895), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n228), .A2(G952), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n604), .A2(new_n609), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n616), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  NAND4_X1  g718(.A1(new_n853), .A2(G210), .A3(new_n858), .A4(G902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n853), .A2(G902), .A3(new_n858), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n853), .A2(new_n910), .A3(new_n858), .A4(G902), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n612), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n904), .A2(new_n906), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n901), .B(new_n907), .C1(new_n912), .C2(new_n913), .ZN(G51));
  INV_X1    g728(.A(new_n786), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n909), .A2(new_n915), .A3(new_n911), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n787), .B(KEYINPUT57), .Z(new_n917));
  AND3_X1   g731(.A1(new_n853), .A2(KEYINPUT54), .A3(new_n858), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n859), .ZN(new_n919));
  AOI22_X1  g733(.A1(KEYINPUT122), .A2(new_n916), .B1(new_n919), .B2(new_n547), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n909), .A2(new_n921), .A3(new_n915), .A4(new_n911), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n901), .B1(new_n920), .B2(new_n922), .ZN(G54));
  AND2_X1   g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n909), .A2(new_n911), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n407), .A3(new_n414), .ZN(new_n926));
  INV_X1    g740(.A(new_n901), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n407), .A2(new_n414), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n909), .A2(new_n928), .A3(new_n911), .A4(new_n924), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(G60));
  OAI21_X1  g744(.A(new_n627), .B1(new_n629), .B2(new_n626), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n852), .A2(new_n860), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT59), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n932), .B(new_n935), .C1(new_n918), .C2(new_n859), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n927), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT60), .Z(new_n941));
  NAND3_X1  g755(.A1(new_n853), .A2(new_n858), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n901), .B1(new_n942), .B2(new_n252), .ZN(new_n943));
  INV_X1    g757(.A(new_n667), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n942), .ZN(new_n945));
  XNOR2_X1  g759(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G66));
  OAI21_X1  g761(.A(G953), .B1(new_n471), .B2(new_n585), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT124), .ZN(new_n949));
  INV_X1    g763(.A(new_n818), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n828), .A2(new_n829), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n949), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n604), .B1(G898), .B2(new_n228), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  NAND2_X1  g769(.A1(new_n325), .A2(new_n327), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n313), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT125), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n681), .A2(new_n710), .A3(new_n750), .ZN(new_n961));
  OR3_X1    g775(.A1(new_n705), .A2(KEYINPUT62), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT62), .B1(new_n705), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n686), .A2(new_n688), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n371), .A2(new_n964), .A3(new_n792), .A4(new_n827), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n809), .B2(new_n811), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(new_n803), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n228), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n801), .B2(new_n802), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n757), .A2(new_n740), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n805), .A2(new_n685), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n771), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n777), .B1(new_n809), .B2(new_n811), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n960), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n968), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n517), .B2(new_n676), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G72));
  XNOR2_X1  g794(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n952), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n974), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n360), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n901), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n967), .B2(new_n984), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n699), .ZN(new_n989));
  INV_X1    g803(.A(new_n983), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n986), .A2(new_n699), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n848), .A2(new_n851), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n987), .A2(new_n989), .A3(KEYINPUT127), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G57));
endmodule


