//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(KEYINPUT78), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n187), .A2(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n195), .B(new_n188), .C1(new_n196), .C2(KEYINPUT23), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n197), .A2(G110), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(KEYINPUT78), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT16), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  OR3_X1    g017(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(G146), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n197), .A2(G110), .ZN(new_n209));
  XOR2_X1   g023(.A(new_n209), .B(KEYINPUT77), .Z(new_n210));
  INV_X1    g024(.A(new_n205), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n202), .B2(new_n204), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n211), .A2(new_n212), .B1(new_n191), .B2(new_n192), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n208), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G137), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n215), .B(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G902), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n208), .B(new_n218), .C1(new_n210), .C2(new_n213), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(KEYINPUT25), .A3(new_n221), .A4(new_n222), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(KEYINPUT79), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(G234), .B2(new_n221), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n230), .A3(new_n224), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n229), .A2(G902), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n222), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n235), .B(KEYINPUT80), .Z(new_n236));
  OAI21_X1  g050(.A(new_n232), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G137), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(G134), .B2(new_n244), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n241), .A2(KEYINPUT11), .A3(G137), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n240), .B(new_n242), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT11), .B1(new_n241), .B2(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n244), .A3(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n240), .B1(new_n251), .B2(new_n242), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n239), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n242), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n247), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT64), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  AOI21_X1  g080(.A(G146), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n206), .A2(G143), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n259), .B(new_n262), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT64), .B(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n206), .A2(G143), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n260), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n268), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n270), .B2(G146), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n259), .B1(new_n276), .B2(new_n262), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n272), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n270), .B2(G146), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G128), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT1), .B1(new_n263), .B2(G146), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n272), .A2(new_n285), .A3(KEYINPUT1), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(G128), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n287), .A2(new_n288), .A3(new_n276), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n287), .B2(new_n276), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n244), .B2(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n244), .A2(G134), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n241), .A2(KEYINPUT67), .A3(G137), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G131), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n247), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n258), .A2(new_n278), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n187), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G113), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT2), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G113), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n313), .A3(KEYINPUT71), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT71), .B1(new_n306), .B2(new_n313), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n313), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT73), .B1(new_n321), .B2(new_n314), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT28), .B1(new_n300), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n291), .A2(new_n299), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n278), .A2(new_n256), .A3(new_n253), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n248), .A2(new_n252), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n264), .A2(new_n266), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n268), .B1(new_n329), .B2(new_n206), .ZN(new_n330));
  INV_X1    g144(.A(new_n262), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT65), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n273), .A3(new_n269), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n333), .B2(KEYINPUT66), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT66), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n335), .A3(new_n273), .A4(new_n269), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n297), .A2(new_n247), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n297), .B2(new_n247), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n334), .A2(new_n336), .B1(new_n291), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n315), .A2(new_n316), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n327), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n324), .B1(new_n343), .B2(KEYINPUT28), .ZN(new_n344));
  INV_X1    g158(.A(G210), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n345), .A2(G237), .A3(G953), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT27), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G101), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n238), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT66), .B1(new_n274), .B2(new_n277), .ZN(new_n353));
  INV_X1    g167(.A(new_n328), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n291), .A2(new_n340), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n342), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT28), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n327), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT74), .A3(new_n349), .ZN(new_n362));
  INV_X1    g176(.A(new_n342), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n355), .A2(new_n356), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n325), .B2(new_n326), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n327), .A3(new_n350), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT31), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n355), .A2(new_n356), .A3(new_n364), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n300), .B2(new_n364), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n352), .B1(new_n372), .B2(new_n363), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT31), .A3(new_n350), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n351), .A2(new_n362), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(G472), .A2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n344), .A2(new_n349), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n287), .A2(new_n276), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT70), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n287), .A2(new_n276), .A3(new_n288), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n298), .B1(new_n384), .B2(new_n282), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n257), .A2(new_n333), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT30), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n342), .B1(new_n387), .B2(new_n371), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n388), .A2(new_n352), .A3(new_n350), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n379), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n349), .A2(new_n379), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n300), .A2(new_n323), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(new_n352), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n360), .B(new_n391), .C1(new_n393), .C2(new_n359), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT76), .ZN(new_n395));
  AOI21_X1  g209(.A(G902), .B1(new_n394), .B2(KEYINPUT76), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n378), .A2(KEYINPUT32), .B1(new_n397), .B2(G472), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n375), .B2(new_n377), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT74), .B1(new_n361), .B2(new_n349), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n238), .B(new_n350), .C1(new_n358), .C2(new_n360), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT31), .B1(new_n373), .B2(new_n350), .ZN(new_n403));
  NOR4_X1   g217(.A1(new_n388), .A2(new_n369), .A3(new_n352), .A4(new_n349), .ZN(new_n404));
  OAI22_X1  g218(.A1(new_n401), .A2(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT75), .A3(new_n376), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n237), .B1(new_n398), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT9), .B(G234), .ZN(new_n410));
  OAI21_X1  g224(.A(G221), .B1(new_n410), .B2(G902), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(KEYINPUT81), .Z(new_n412));
  INV_X1    g226(.A(G104), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT3), .B1(new_n413), .B2(G107), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G104), .ZN(new_n417));
  INV_X1    g231(.A(G101), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(G107), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n414), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n413), .A2(G107), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n416), .A2(G104), .ZN(new_n422));
  OAI21_X1  g236(.A(G101), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n291), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n424), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT1), .B1(new_n270), .B2(G146), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n280), .B1(G128), .B2(new_n429), .ZN(new_n430));
  AND4_X1   g244(.A1(new_n281), .A2(new_n271), .A3(G128), .A4(new_n272), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n414), .A2(new_n417), .A3(new_n419), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G101), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(G101), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT4), .A3(new_n420), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n278), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n427), .A2(new_n433), .A3(new_n439), .A4(new_n257), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT82), .ZN(new_n442));
  INV_X1    g256(.A(G227), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n442), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n440), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n282), .B(new_n424), .C1(new_n289), .C2(new_n290), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n432), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n354), .A2(KEYINPUT12), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n257), .B1(new_n450), .B2(new_n432), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n453), .B1(KEYINPUT12), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n445), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n433), .A2(new_n439), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n257), .B1(new_n458), .B2(new_n427), .ZN(new_n459));
  INV_X1    g273(.A(new_n440), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n459), .A2(new_n446), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n445), .B1(new_n455), .B2(new_n440), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G469), .B1(new_n467), .B2(G902), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n412), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G214), .B1(G237), .B2(G902), .ZN(new_n470));
  NAND2_X1  g284(.A1(G234), .A2(G237), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n471), .A2(G902), .A3(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(G898), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n471), .A2(G952), .A3(new_n216), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n333), .A2(G125), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n203), .B(new_n282), .C1(new_n289), .C2(new_n290), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n216), .A2(G224), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT7), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n312), .A2(KEYINPUT5), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(G113), .C1(KEYINPUT5), .C2(new_n301), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n313), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n420), .A2(new_n423), .A3(KEYINPUT85), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT8), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n479), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n495), .B2(new_n481), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT86), .B(new_n482), .C1(new_n478), .C2(new_n479), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n428), .A2(new_n485), .A3(new_n313), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n438), .A2(new_n436), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n490), .B(new_n501), .C1(new_n342), .C2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n493), .B(KEYINPUT87), .C1(new_n496), .C2(new_n497), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n501), .B1(new_n342), .B2(new_n502), .ZN(new_n506));
  INV_X1    g320(.A(new_n490), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(KEYINPUT84), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n508), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n495), .B(new_n480), .Z(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G210), .B1(G237), .B2(G902), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n505), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n505), .B2(new_n514), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n470), .B(new_n477), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n521));
  INV_X1    g335(.A(G214), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n522), .A2(G237), .A3(G953), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G143), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n329), .B2(new_n523), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n525), .B2(G131), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n521), .A3(G131), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT17), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n211), .A2(new_n212), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n525), .A2(new_n521), .A3(G131), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n531), .A2(new_n526), .B1(G131), .B2(new_n525), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n529), .B(new_n530), .C1(new_n532), .C2(KEYINPUT17), .ZN(new_n533));
  XNOR2_X1  g347(.A(G113), .B(G122), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(new_n413), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n201), .B(new_n206), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n240), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n525), .A2(G131), .ZN(new_n539));
  OAI221_X1 g353(.A(new_n536), .B1(new_n525), .B2(new_n538), .C1(new_n539), .C2(new_n537), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(KEYINPUT19), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n201), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n201), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n205), .B1(new_n546), .B2(G146), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(KEYINPUT90), .B(new_n205), .C1(new_n546), .C2(G146), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n532), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n535), .B1(new_n551), .B2(new_n540), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n520), .B1(new_n541), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n552), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n520), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n535), .B1(new_n533), .B2(new_n540), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n221), .B1(new_n541), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n554), .A2(new_n559), .B1(G475), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n270), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n189), .A2(G143), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G134), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n302), .A2(G122), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n416), .B1(new_n567), .B2(KEYINPUT14), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n302), .A2(G122), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n570), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n410), .A2(new_n228), .A3(G953), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n329), .A2(new_n189), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n241), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n576), .B2(new_n565), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n580));
  INV_X1    g394(.A(new_n565), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT13), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n582), .B2(new_n577), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n241), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n567), .A2(new_n569), .A3(G107), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n570), .A2(new_n416), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n573), .B(new_n574), .C1(new_n584), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n574), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n580), .A3(new_n577), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n562), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n519), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n409), .A2(new_n469), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NOR3_X1   g417(.A1(new_n375), .A2(new_n399), .A3(new_n377), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT75), .B1(new_n405), .B2(new_n376), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT92), .B1(new_n375), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n405), .A2(new_n608), .A3(new_n221), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G472), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n237), .ZN(new_n611));
  AND4_X1   g425(.A1(new_n606), .A2(new_n610), .A3(new_n611), .A4(new_n469), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT93), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n589), .A2(new_n595), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT33), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n589), .A2(new_n595), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(G478), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n597), .A2(new_n221), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n596), .B2(new_n597), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n562), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n519), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G104), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n629));
  INV_X1    g443(.A(new_n599), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n562), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n519), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n470), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n505), .A2(new_n514), .ZN(new_n634));
  INV_X1    g448(.A(new_n515), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n633), .B1(new_n636), .B2(new_n516), .ZN(new_n637));
  INV_X1    g451(.A(new_n631), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(KEYINPUT95), .A3(new_n477), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n613), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  XNOR2_X1  g457(.A(new_n214), .B(KEYINPUT96), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n219), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n232), .B1(new_n234), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n232), .B(KEYINPUT97), .C1(new_n234), .C2(new_n646), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n469), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n601), .A3(new_n606), .A4(new_n610), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n398), .A2(new_n408), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n470), .B1(new_n517), .B2(new_n518), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n475), .B1(new_n472), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n630), .A2(new_n562), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT98), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n661), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n637), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n656), .A2(new_n652), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NAND2_X1  g481(.A1(new_n636), .A2(new_n516), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n647), .A2(new_n562), .A3(new_n633), .A4(new_n599), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n659), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n469), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n378), .A2(KEYINPUT32), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n350), .B1(new_n388), .B2(new_n352), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n393), .A2(new_n349), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n221), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G472), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n408), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n671), .A2(new_n674), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n329), .ZN(G45));
  AND2_X1   g496(.A1(new_n618), .A2(new_n620), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n561), .A2(G475), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n558), .B1(new_n557), .B2(new_n520), .ZN(new_n685));
  INV_X1    g499(.A(new_n520), .ZN(new_n686));
  AOI211_X1 g500(.A(KEYINPUT20), .B(new_n686), .C1(new_n555), .C2(new_n556), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n688), .A3(new_n660), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n657), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n656), .A2(new_n652), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  INV_X1    g506(.A(new_n411), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT99), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n462), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n462), .B2(new_n694), .ZN(new_n697));
  OAI211_X1 g511(.A(KEYINPUT100), .B(new_n464), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n462), .A2(new_n694), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(new_n700), .A3(G469), .A4(new_n695), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n693), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n409), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n624), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n640), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  AOI211_X1 g522(.A(new_n693), .B(new_n657), .C1(new_n698), .C2(new_n701), .ZN(new_n709));
  INV_X1    g523(.A(new_n600), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n649), .A3(new_n650), .A4(new_n477), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n398), .B2(new_n408), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  INV_X1    g528(.A(G472), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n405), .B2(new_n221), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n370), .A2(new_n374), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n360), .B1(new_n393), .B2(new_n359), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n349), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n377), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n720), .A3(new_n237), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n562), .B2(new_n599), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n630), .A2(KEYINPUT101), .A3(new_n688), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n519), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n702), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n622), .A2(new_n729), .A3(new_n660), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n689), .A2(KEYINPUT102), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n647), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n716), .A2(new_n733), .A3(new_n720), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n702), .A2(new_n732), .A3(new_n637), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  AOI211_X1 g550(.A(G469), .B(G902), .C1(new_n456), .C2(new_n461), .ZN(new_n737));
  NAND2_X1  g551(.A1(G469), .A2(G902), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT103), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n455), .A2(new_n440), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n457), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n433), .A2(new_n439), .ZN(new_n742));
  INV_X1    g556(.A(new_n427), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n258), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n445), .A3(new_n440), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n739), .B1(new_n746), .B2(new_n463), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT104), .B1(new_n737), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  INV_X1    g563(.A(new_n739), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n467), .B2(G469), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n464), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n693), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n636), .A2(new_n470), .A3(new_n516), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n636), .A2(new_n516), .A3(KEYINPUT105), .A4(new_n470), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n732), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n398), .B1(KEYINPUT32), .B2(new_n378), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n611), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n409), .A2(new_n758), .A3(new_n732), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND3_X1  g584(.A1(new_n409), .A2(new_n758), .A3(new_n663), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n683), .A2(new_n562), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT43), .Z(new_n774));
  NAND2_X1  g588(.A1(new_n606), .A2(new_n610), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT108), .B1(new_n775), .B2(new_n647), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n777), .B(new_n733), .C1(new_n606), .C2(new_n610), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(KEYINPUT44), .B(new_n774), .C1(new_n776), .C2(new_n778), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n741), .A2(KEYINPUT45), .A3(new_n745), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n465), .B2(new_n466), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n785), .A3(G469), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n783), .A2(new_n785), .A3(KEYINPUT107), .A4(G469), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n750), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n464), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n792), .B(new_n750), .C1(new_n788), .C2(new_n789), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n411), .B(new_n672), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n756), .A2(new_n757), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n781), .A2(new_n782), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  INV_X1    g612(.A(new_n795), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n611), .A2(new_n689), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(new_n408), .A3(new_n398), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n411), .B1(new_n791), .B2(new_n793), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT47), .B(new_n411), .C1(new_n791), .C2(new_n793), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(G140), .Z(G42));
  NAND2_X1  g621(.A1(new_n698), .A2(new_n701), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT109), .Z(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT110), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n812));
  INV_X1    g626(.A(new_n412), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n611), .A2(new_n813), .A3(new_n470), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n680), .A2(new_n669), .A3(new_n773), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n774), .A2(new_n475), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n702), .A3(new_n799), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT116), .Z(new_n819));
  OAI21_X1  g633(.A(G472), .B1(new_n375), .B2(G902), .ZN(new_n820));
  INV_X1    g634(.A(new_n720), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n647), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n817), .A2(new_n721), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n795), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n809), .A2(new_n813), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n804), .A2(new_n805), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n680), .A2(new_n237), .A3(new_n476), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n799), .A2(new_n702), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n829), .A2(new_n688), .A3(new_n683), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n633), .B1(KEYINPUT115), .B2(KEYINPUT50), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n669), .A2(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n702), .A2(new_n817), .A3(new_n721), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n823), .A2(new_n828), .A3(new_n832), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  INV_X1    g655(.A(new_n709), .ZN(new_n842));
  OAI211_X1 g656(.A(G952), .B(new_n216), .C1(new_n824), .C2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n829), .A2(new_n623), .A3(new_n830), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n819), .A2(new_n761), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n840), .A2(new_n841), .A3(new_n850), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n623), .A2(KEYINPUT111), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n638), .B1(new_n623), .B2(KEYINPUT111), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n519), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n612), .A2(new_n854), .B1(new_n709), .B2(new_n712), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n727), .A2(new_n653), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n409), .B(new_n702), .C1(new_n640), .C2(new_n624), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n602), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n651), .B1(new_n398), .B2(new_n408), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n799), .A3(new_n710), .A4(new_n660), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n730), .A2(new_n731), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n822), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n758), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n771), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n769), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n662), .A2(new_n665), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n859), .A2(new_n867), .B1(new_n709), .B2(new_n862), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n733), .A2(new_n411), .A3(new_n660), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n752), .B2(new_n748), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n725), .A2(new_n657), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n680), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(new_n869), .A3(new_n691), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n666), .A2(new_n873), .A3(new_n691), .A4(new_n735), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT112), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT112), .B1(new_n874), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n874), .A2(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n865), .A3(new_n769), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n882));
  AOI22_X1  g696(.A1(new_n866), .A2(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n768), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n762), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n860), .A2(new_n771), .A3(new_n863), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n602), .A2(new_n653), .A3(new_n727), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n855), .A4(new_n857), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n879), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n881), .A2(new_n882), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n885), .B(KEYINPUT114), .C1(new_n895), .C2(new_n884), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n885), .A2(KEYINPUT114), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n851), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n816), .B1(new_n898), .B2(new_n899), .ZN(G75));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n866), .A2(new_n879), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n881), .A2(new_n882), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n221), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT56), .B1(new_n904), .B2(G210), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n512), .B(new_n513), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n901), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n883), .A2(new_n345), .A3(new_n221), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT118), .B(new_n907), .C1(new_n910), .C2(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n216), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n904), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT119), .B1(new_n883), .B2(new_n221), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n635), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n912), .A2(new_n919), .ZN(G51));
  NAND2_X1  g734(.A1(new_n456), .A2(new_n461), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n883), .B(KEYINPUT54), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n739), .B(KEYINPUT57), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n915), .A2(new_n916), .A3(new_n788), .A4(new_n789), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n913), .B1(new_n924), .B2(new_n925), .ZN(G54));
  NAND2_X1  g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT120), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n915), .A2(new_n916), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n556), .A3(new_n555), .ZN(new_n930));
  INV_X1    g744(.A(new_n913), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n915), .A2(new_n916), .A3(new_n557), .A4(new_n928), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G60));
  AND2_X1   g747(.A1(new_n615), .A2(new_n617), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(new_n619), .Z(new_n936));
  OR2_X1    g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n922), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n936), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n897), .A2(new_n896), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n934), .B2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n769), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n945), .A2(new_n877), .A3(new_n878), .ZN(new_n946));
  INV_X1    g760(.A(new_n882), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n892), .B2(new_n880), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n913), .B1(new_n949), .B2(new_n236), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n644), .B(new_n645), .Z(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n944), .C1(new_n946), .C2(new_n948), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT61), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n236), .B1(new_n883), .B2(new_n943), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(new_n953), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT123), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n931), .A3(new_n953), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n959), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(G66));
  INV_X1    g778(.A(G224), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n473), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n858), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(G953), .ZN(new_n968));
  INV_X1    g782(.A(G898), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n512), .B1(new_n969), .B2(G953), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n968), .B(new_n970), .Z(G69));
  XNOR2_X1  g785(.A(new_n372), .B(new_n546), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n216), .A2(G900), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n666), .A2(new_n691), .A3(new_n735), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n666), .A2(new_n691), .A3(new_n735), .A4(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n760), .A2(new_n611), .A3(new_n872), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n771), .B1(new_n980), .B2(new_n794), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n806), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n797), .A2(new_n769), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n974), .B1(new_n983), .B2(new_n216), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n973), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI211_X1 g800(.A(KEYINPUT126), .B(new_n974), .C1(new_n983), .C2(new_n216), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n979), .A2(new_n988), .A3(new_n681), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n681), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n977), .B2(new_n978), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(KEYINPUT125), .A3(new_n988), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n673), .B1(new_n852), .B2(new_n853), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n799), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n806), .B1(new_n409), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n797), .B(new_n998), .C1(new_n993), .C2(new_n988), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  OAI22_X1  g815(.A1(new_n986), .A2(new_n987), .B1(new_n1001), .B2(new_n973), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1003));
  OAI21_X1  g817(.A(G953), .B1(new_n443), .B2(new_n658), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n999), .B1(new_n991), .B2(new_n994), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n972), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1006), .B(new_n1007), .C1(new_n987), .C2(new_n986), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1003), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1004), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n983), .B2(new_n858), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n913), .B1(new_n1014), .B2(new_n389), .ZN(new_n1015));
  INV_X1    g829(.A(new_n389), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n676), .A3(new_n1013), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1015), .B1(new_n895), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1005), .A2(new_n967), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n676), .B1(new_n1019), .B2(new_n1013), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1018), .A2(new_n1020), .ZN(G57));
endmodule


