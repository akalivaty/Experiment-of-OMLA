

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n724) );
  NOR2_X1 U558 ( .A1(n740), .A2(G168), .ZN(n742) );
  NAND2_X1 U559 ( .A1(n758), .A2(G286), .ZN(n747) );
  OR2_X1 U560 ( .A1(n734), .A2(n733), .ZN(n523) );
  AND2_X1 U561 ( .A1(n933), .A2(n834), .ZN(n524) );
  NAND2_X1 U562 ( .A1(n788), .A2(n787), .ZN(n525) );
  XNOR2_X1 U563 ( .A(KEYINPUT31), .B(n746), .ZN(n526) );
  XNOR2_X1 U564 ( .A(n700), .B(KEYINPUT94), .ZN(n701) );
  XNOR2_X1 U565 ( .A(n702), .B(n701), .ZN(n704) );
  INV_X1 U566 ( .A(n748), .ZN(n730) );
  INV_X1 U567 ( .A(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U568 ( .A1(n523), .A2(n526), .ZN(n758) );
  NOR2_X1 U569 ( .A1(n748), .A2(G2084), .ZN(n735) );
  NAND2_X1 U570 ( .A1(n699), .A2(n800), .ZN(n748) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n542) );
  NOR2_X1 U572 ( .A1(n821), .A2(n524), .ZN(n822) );
  NOR2_X1 U573 ( .A1(G2105), .A2(n549), .ZN(n895) );
  NOR2_X1 U574 ( .A1(G651), .A2(n645), .ZN(n664) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n655) );
  NAND2_X1 U576 ( .A1(G89), .A2(n655), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT4), .B(n527), .Z(n528) );
  XNOR2_X1 U578 ( .A(n528), .B(KEYINPUT73), .ZN(n532) );
  INV_X1 U579 ( .A(G651), .ZN(n534) );
  XNOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .ZN(n529) );
  XOR2_X1 U581 ( .A(n529), .B(KEYINPUT66), .Z(n645) );
  OR2_X1 U582 ( .A1(n534), .A2(n645), .ZN(n530) );
  XNOR2_X1 U583 ( .A(KEYINPUT67), .B(n530), .ZN(n659) );
  NAND2_X1 U584 ( .A1(G76), .A2(n659), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n533), .B(KEYINPUT5), .ZN(n540) );
  NAND2_X1 U587 ( .A1(G51), .A2(n664), .ZN(n537) );
  NOR2_X1 U588 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n535), .Z(n656) );
  NAND2_X1 U590 ( .A1(G63), .A2(n656), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U594 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U595 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X2 U596 ( .A(KEYINPUT17), .B(n542), .Z(n894) );
  NAND2_X1 U597 ( .A1(G137), .A2(n894), .ZN(n545) );
  INV_X1 U598 ( .A(G2104), .ZN(n549) );
  AND2_X1 U599 ( .A1(G2105), .A2(G2104), .ZN(n900) );
  NAND2_X1 U600 ( .A1(n900), .A2(G113), .ZN(n543) );
  XNOR2_X1 U601 ( .A(n543), .B(KEYINPUT64), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT65), .ZN(n548) );
  AND2_X1 U604 ( .A1(n549), .A2(G2105), .ZN(n898) );
  NAND2_X1 U605 ( .A1(G125), .A2(n898), .ZN(n547) );
  AND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n698) );
  NAND2_X1 U607 ( .A1(G101), .A2(n895), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(n550), .Z(n696) );
  AND2_X1 U609 ( .A1(n698), .A2(n696), .ZN(G160) );
  XNOR2_X1 U610 ( .A(G2451), .B(G2446), .ZN(n560) );
  XOR2_X1 U611 ( .A(G2430), .B(KEYINPUT105), .Z(n552) );
  XNOR2_X1 U612 ( .A(G2454), .B(G2435), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n552), .B(n551), .ZN(n556) );
  XOR2_X1 U614 ( .A(G2438), .B(KEYINPUT104), .Z(n554) );
  XNOR2_X1 U615 ( .A(G1341), .B(G1348), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U617 ( .A(n556), .B(n555), .Z(n558) );
  XNOR2_X1 U618 ( .A(G2443), .B(G2427), .ZN(n557) );
  XNOR2_X1 U619 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n560), .B(n559), .ZN(n561) );
  AND2_X1 U621 ( .A1(n561), .A2(G14), .ZN(G401) );
  NAND2_X1 U622 ( .A1(G52), .A2(n664), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G64), .A2(n656), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G90), .A2(n655), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G77), .A2(n659), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n566), .Z(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(G171) );
  INV_X1 U630 ( .A(G171), .ZN(G301) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  INV_X1 U632 ( .A(G82), .ZN(G220) );
  NAND2_X1 U633 ( .A1(G88), .A2(n655), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G75), .A2(n659), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G50), .A2(n664), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G62), .A2(n656), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(G166) );
  NAND2_X1 U640 ( .A1(G138), .A2(n894), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G102), .A2(n895), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G126), .A2(n898), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G114), .A2(n900), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(G164) );
  NAND2_X1 U647 ( .A1(G94), .A2(G452), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT69), .ZN(G173) );
  XOR2_X1 U649 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n583) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n583), .B(n582), .ZN(G223) );
  XOR2_X1 U652 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n585) );
  INV_X1 U653 ( .A(G223), .ZN(n839) );
  NAND2_X1 U654 ( .A1(G567), .A2(n839), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n585), .B(n584), .ZN(G234) );
  NAND2_X1 U656 ( .A1(G56), .A2(n656), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT14), .B(n586), .Z(n592) );
  NAND2_X1 U658 ( .A1(n655), .A2(G81), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G68), .A2(n659), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n664), .A2(G43), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n1014) );
  INV_X1 U666 ( .A(G860), .ZN(n614) );
  OR2_X1 U667 ( .A1(n1014), .A2(n614), .ZN(G153) );
  NAND2_X1 U668 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G54), .A2(n664), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G66), .A2(n656), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G92), .A2(n655), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G79), .A2(n659), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT15), .ZN(n998) );
  INV_X1 U677 ( .A(G868), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n998), .A2(n610), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U680 ( .A1(G53), .A2(n664), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G65), .A2(n656), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G91), .A2(n655), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G78), .A2(n659), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n1006) );
  INV_X1 U687 ( .A(n1006), .ZN(G299) );
  NOR2_X1 U688 ( .A1(G286), .A2(n610), .ZN(n611) );
  XNOR2_X1 U689 ( .A(n611), .B(KEYINPUT74), .ZN(n613) );
  NOR2_X1 U690 ( .A1(G299), .A2(G868), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n614), .A2(G559), .ZN(n615) );
  INV_X1 U693 ( .A(n998), .ZN(n631) );
  NAND2_X1 U694 ( .A1(n615), .A2(n631), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U696 ( .A1(G868), .A2(n1014), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT75), .B(n617), .Z(n620) );
  NAND2_X1 U698 ( .A1(G868), .A2(n631), .ZN(n618) );
  NOR2_X1 U699 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U701 ( .A(KEYINPUT76), .B(n621), .ZN(G282) );
  XNOR2_X1 U702 ( .A(G2100), .B(KEYINPUT77), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n898), .A2(G123), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n622), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G111), .A2(n900), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G135), .A2(n894), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G99), .A2(n895), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n932) );
  XNOR2_X1 U711 ( .A(n932), .B(G2096), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U713 ( .A1(n631), .A2(G559), .ZN(n676) );
  XNOR2_X1 U714 ( .A(n1014), .B(n676), .ZN(n632) );
  NOR2_X1 U715 ( .A1(n632), .A2(G860), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G93), .A2(n655), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G80), .A2(n659), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U719 ( .A(KEYINPUT78), .B(n635), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G55), .A2(n664), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G67), .A2(n656), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n673) );
  XNOR2_X1 U724 ( .A(n640), .B(n673), .ZN(G145) );
  NAND2_X1 U725 ( .A1(G49), .A2(n664), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U728 ( .A1(n656), .A2(n643), .ZN(n644) );
  XOR2_X1 U729 ( .A(KEYINPUT79), .B(n644), .Z(n647) );
  NAND2_X1 U730 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U732 ( .A1(n659), .A2(G72), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n655), .A2(G85), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U735 ( .A1(G47), .A2(n664), .ZN(n650) );
  XOR2_X1 U736 ( .A(KEYINPUT68), .B(n650), .Z(n651) );
  NOR2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n656), .A2(G60), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(G290) );
  NAND2_X1 U740 ( .A1(G86), .A2(n655), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G61), .A2(n656), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n659), .A2(G73), .ZN(n660) );
  XOR2_X1 U744 ( .A(KEYINPUT2), .B(n660), .Z(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n663), .B(KEYINPUT80), .ZN(n666) );
  NAND2_X1 U747 ( .A1(G48), .A2(n664), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n666), .A2(n665), .ZN(G305) );
  NOR2_X1 U749 ( .A1(G868), .A2(n673), .ZN(n667) );
  XOR2_X1 U750 ( .A(n667), .B(KEYINPUT82), .Z(n679) );
  XNOR2_X1 U751 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n669) );
  XNOR2_X1 U752 ( .A(G288), .B(G166), .ZN(n668) );
  XNOR2_X1 U753 ( .A(n669), .B(n668), .ZN(n672) );
  XNOR2_X1 U754 ( .A(n1006), .B(G290), .ZN(n670) );
  XNOR2_X1 U755 ( .A(n670), .B(n1014), .ZN(n671) );
  XNOR2_X1 U756 ( .A(n672), .B(n671), .ZN(n675) );
  XNOR2_X1 U757 ( .A(G305), .B(n673), .ZN(n674) );
  XNOR2_X1 U758 ( .A(n675), .B(n674), .ZN(n911) );
  XOR2_X1 U759 ( .A(n911), .B(n676), .Z(n677) );
  NAND2_X1 U760 ( .A1(G868), .A2(n677), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XNOR2_X1 U763 ( .A(n680), .B(KEYINPUT83), .ZN(n681) );
  XNOR2_X1 U764 ( .A(n681), .B(KEYINPUT20), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n682), .A2(G2090), .ZN(n683) );
  XNOR2_X1 U766 ( .A(n683), .B(KEYINPUT21), .ZN(n684) );
  XNOR2_X1 U767 ( .A(n684), .B(KEYINPUT84), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XOR2_X1 U769 ( .A(KEYINPUT85), .B(G44), .Z(n686) );
  XNOR2_X1 U770 ( .A(KEYINPUT3), .B(n686), .ZN(G218) );
  XOR2_X1 U771 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U772 ( .A1(G219), .A2(G220), .ZN(n687) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U774 ( .A1(G218), .A2(n688), .ZN(n689) );
  NAND2_X1 U775 ( .A1(G96), .A2(n689), .ZN(n844) );
  AND2_X1 U776 ( .A1(G2106), .A2(n844), .ZN(n694) );
  NAND2_X1 U777 ( .A1(G69), .A2(G120), .ZN(n690) );
  NOR2_X1 U778 ( .A1(G237), .A2(n690), .ZN(n691) );
  NAND2_X1 U779 ( .A1(G108), .A2(n691), .ZN(n843) );
  NAND2_X1 U780 ( .A1(G567), .A2(n843), .ZN(n692) );
  XOR2_X1 U781 ( .A(KEYINPUT86), .B(n692), .Z(n693) );
  NOR2_X1 U782 ( .A1(n694), .A2(n693), .ZN(G319) );
  INV_X1 U783 ( .A(G319), .ZN(n919) );
  NAND2_X1 U784 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U785 ( .A1(n919), .A2(n695), .ZN(n842) );
  NAND2_X1 U786 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U787 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U788 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n729) );
  AND2_X1 U789 ( .A1(G40), .A2(n696), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n799) );
  INV_X1 U791 ( .A(n799), .ZN(n699) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n800) );
  NAND2_X1 U793 ( .A1(G2072), .A2(n730), .ZN(n702) );
  XOR2_X1 U794 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n700) );
  AND2_X1 U795 ( .A1(G1956), .A2(n748), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n723) );
  NAND2_X1 U797 ( .A1(n1006), .A2(n723), .ZN(n722) );
  INV_X1 U798 ( .A(G1341), .ZN(n981) );
  NOR2_X1 U799 ( .A1(n730), .A2(n981), .ZN(n705) );
  NAND2_X1 U800 ( .A1(KEYINPUT26), .A2(n705), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n707), .A2(KEYINPUT95), .ZN(n712) );
  INV_X1 U802 ( .A(KEYINPUT95), .ZN(n710) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n730), .ZN(n706) );
  XNOR2_X1 U804 ( .A(KEYINPUT26), .B(n706), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n1014), .A2(n713), .ZN(n717) );
  NAND2_X1 U809 ( .A1(G1348), .A2(n748), .ZN(n715) );
  NAND2_X1 U810 ( .A1(G2067), .A2(n730), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n998), .A2(n718), .ZN(n716) );
  OR2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n998), .A2(n718), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n727) );
  NOR2_X1 U817 ( .A1(n1006), .A2(n723), .ZN(n725) );
  XNOR2_X1 U818 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n729), .B(n728), .ZN(n734) );
  NOR2_X1 U821 ( .A1(n730), .A2(G1961), .ZN(n732) );
  XOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .Z(n960) );
  NOR2_X1 U823 ( .A1(n748), .A2(n960), .ZN(n731) );
  NOR2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n743) );
  NOR2_X1 U825 ( .A1(n743), .A2(G301), .ZN(n733) );
  XNOR2_X1 U826 ( .A(KEYINPUT97), .B(KEYINPUT30), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G8), .A2(n748), .ZN(n783) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n783), .ZN(n760) );
  XNOR2_X1 U829 ( .A(n735), .B(KEYINPUT92), .ZN(n757) );
  INV_X1 U830 ( .A(n757), .ZN(n736) );
  NAND2_X1 U831 ( .A1(n736), .A2(G8), .ZN(n737) );
  NOR2_X1 U832 ( .A1(n760), .A2(n737), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U834 ( .A(n742), .B(n741), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n743), .A2(G301), .ZN(n744) );
  NAND2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U837 ( .A(KEYINPUT99), .B(n747), .Z(n753) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n783), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n748), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U841 ( .A1(G303), .A2(n751), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n754), .A2(G8), .ZN(n756) );
  XNOR2_X1 U844 ( .A(KEYINPUT100), .B(KEYINPUT32), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n756), .B(n755), .ZN(n764) );
  NAND2_X1 U846 ( .A1(n757), .A2(G8), .ZN(n762) );
  INV_X1 U847 ( .A(n758), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n779) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n1009) );
  NOR2_X1 U853 ( .A1(n765), .A2(n1009), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n779), .A2(n766), .ZN(n767) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  NAND2_X1 U856 ( .A1(n767), .A2(n1007), .ZN(n773) );
  NAND2_X1 U857 ( .A1(n1009), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n768), .A2(n783), .ZN(n770) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n1003) );
  INV_X1 U860 ( .A(n1003), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n774) );
  INV_X1 U862 ( .A(n774), .ZN(n771) );
  OR2_X1 U863 ( .A1(n783), .A2(n771), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n776) );
  AND2_X1 U865 ( .A1(n774), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n788) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  AND2_X1 U870 ( .A1(n780), .A2(n783), .ZN(n786) );
  NOR2_X1 U871 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XOR2_X1 U872 ( .A(n781), .B(KEYINPUT24), .Z(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT91), .B(n784), .Z(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G140), .A2(n894), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G104), .A2(n895), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n791), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G128), .A2(n898), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G116), .A2(n900), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT35), .B(n794), .Z(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT88), .B(n795), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n798), .ZN(n907) );
  XNOR2_X1 U887 ( .A(KEYINPUT37), .B(G2067), .ZN(n832) );
  NOR2_X1 U888 ( .A1(n907), .A2(n832), .ZN(n929) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n834) );
  NAND2_X1 U890 ( .A1(n929), .A2(n834), .ZN(n801) );
  XOR2_X1 U891 ( .A(KEYINPUT89), .B(n801), .Z(n830) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n824) );
  INV_X1 U893 ( .A(n824), .ZN(n1012) );
  NAND2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n1001) );
  NAND2_X1 U895 ( .A1(n1012), .A2(n1001), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n802), .A2(n834), .ZN(n803) );
  XOR2_X1 U897 ( .A(KEYINPUT87), .B(n803), .Z(n804) );
  NAND2_X1 U898 ( .A1(n830), .A2(n804), .ZN(n821) );
  NAND2_X1 U899 ( .A1(G95), .A2(n895), .ZN(n806) );
  NAND2_X1 U900 ( .A1(G107), .A2(n900), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n894), .A2(G131), .ZN(n807) );
  XOR2_X1 U903 ( .A(KEYINPUT90), .B(n807), .Z(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n898), .A2(G119), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n889) );
  NAND2_X1 U907 ( .A1(G1991), .A2(n889), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G141), .A2(n894), .ZN(n813) );
  NAND2_X1 U909 ( .A1(G129), .A2(n898), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n895), .A2(G105), .ZN(n814) );
  XOR2_X1 U912 ( .A(KEYINPUT38), .B(n814), .Z(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n900), .A2(G117), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n877) );
  NAND2_X1 U916 ( .A1(G1996), .A2(n877), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n933) );
  NAND2_X1 U918 ( .A1(n525), .A2(n822), .ZN(n837) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n877), .ZN(n823) );
  XOR2_X1 U920 ( .A(KEYINPUT101), .B(n823), .Z(n924) );
  NOR2_X1 U921 ( .A1(G1991), .A2(n889), .ZN(n934) );
  NOR2_X1 U922 ( .A1(n934), .A2(n824), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n825), .B(KEYINPUT102), .ZN(n826) );
  NOR2_X1 U924 ( .A1(n933), .A2(n826), .ZN(n827) );
  NOR2_X1 U925 ( .A1(n924), .A2(n827), .ZN(n828) );
  XOR2_X1 U926 ( .A(n828), .B(KEYINPUT39), .Z(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT103), .B(n829), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U929 ( .A1(n907), .A2(n832), .ZN(n928) );
  NAND2_X1 U930 ( .A1(n833), .A2(n928), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(KEYINPUT40), .B(n838), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U936 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G69), .ZN(G235) );
  NOR2_X1 U943 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  XOR2_X1 U945 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n846) );
  XNOR2_X1 U946 ( .A(KEYINPUT106), .B(G2678), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2072), .Z(n848) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2090), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2100), .B(G2096), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U954 ( .A(G2078), .B(G2084), .Z(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1966), .B(G1981), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n866) );
  XOR2_X1 U959 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U960 ( .A(G1961), .B(KEYINPUT109), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U962 ( .A(G1956), .B(G1971), .Z(n860) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1976), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(G2474), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U969 ( .A1(G124), .A2(n898), .ZN(n867) );
  XOR2_X1 U970 ( .A(KEYINPUT44), .B(n867), .Z(n868) );
  XNOR2_X1 U971 ( .A(n868), .B(KEYINPUT111), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G136), .A2(n894), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G100), .A2(n895), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G112), .A2(n900), .ZN(n871) );
  NAND2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT112), .B(n875), .ZN(G162) );
  XOR2_X1 U979 ( .A(G160), .B(n932), .Z(n876) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(n893) );
  XOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n888) );
  NAND2_X1 U982 ( .A1(G130), .A2(n898), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G118), .A2(n900), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G142), .A2(n894), .ZN(n881) );
  NAND2_X1 U986 ( .A1(G106), .A2(n895), .ZN(n880) );
  NAND2_X1 U987 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U988 ( .A(KEYINPUT113), .B(n882), .ZN(n883) );
  XNOR2_X1 U989 ( .A(KEYINPUT45), .B(n883), .ZN(n884) );
  NOR2_X1 U990 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U991 ( .A(G164), .B(n886), .ZN(n887) );
  XNOR2_X1 U992 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n891), .B(G162), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n909) );
  NAND2_X1 U996 ( .A1(G139), .A2(n894), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G103), .A2(n895), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n898), .A2(G127), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n899), .B(KEYINPUT114), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n900), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n903), .Z(n904) );
  NOR2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(KEYINPUT115), .B(n906), .Z(n937) );
  XNOR2_X1 U1006 ( .A(n907), .B(n937), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(n911), .B(G301), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n912), .B(n998), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n913), .B(G286), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(KEYINPUT49), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n916), .B(KEYINPUT117), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n920), .B(KEYINPUT116), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1023 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n927) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(KEYINPUT51), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n927), .B(n926), .ZN(n946) );
  INV_X1 U1028 ( .A(n928), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n944) );
  XOR2_X1 U1030 ( .A(G2084), .B(G160), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1034 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1045 ( .A(G2084), .B(G34), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT54), .ZN(n970) );
  XNOR2_X1 U1047 ( .A(G2090), .B(G35), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n952), .B(KEYINPUT120), .ZN(n967) );
  XOR2_X1 U1049 ( .A(G1991), .B(G25), .Z(n953) );
  NAND2_X1 U1050 ( .A1(G28), .A2(n953), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(KEYINPUT121), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(G2072), .B(G33), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G1996), .B(G32), .Z(n962) );
  XOR2_X1 U1057 ( .A(G27), .B(KEYINPUT122), .Z(n959) );
  XNOR2_X1 U1058 ( .A(n960), .B(n959), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n965), .B(KEYINPUT53), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT123), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1065 ( .A(KEYINPUT55), .B(n971), .Z(n972) );
  NOR2_X1 U1066 ( .A1(G29), .A2(n972), .ZN(n1028) );
  XOR2_X1 U1067 ( .A(G1966), .B(G21), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G1976), .B(G23), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G22), .B(G1971), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT126), .B(n975), .Z(n977) );
  XNOR2_X1 U1072 ( .A(G1986), .B(G24), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n993) );
  XOR2_X1 U1076 ( .A(G1961), .B(G5), .Z(n991) );
  XNOR2_X1 U1077 ( .A(G19), .B(n981), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G1981), .B(G6), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(G1956), .B(G20), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1082 ( .A(KEYINPUT59), .B(G1348), .Z(n986) );
  XNOR2_X1 U1083 ( .A(G4), .B(n986), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(n989), .B(KEYINPUT60), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1088 ( .A(KEYINPUT61), .B(n994), .Z(n995) );
  NOR2_X1 U1089 ( .A1(G16), .A2(n995), .ZN(n1025) );
  XOR2_X1 U1090 ( .A(G16), .B(KEYINPUT56), .Z(n1023) );
  XNOR2_X1 U1091 ( .A(G171), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1092 ( .A(G166), .B(G1971), .ZN(n996) );
  NAND2_X1 U1093 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n998), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1021) );
  XNOR2_X1 U1097 ( .A(G168), .B(G1966), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(n1005), .B(KEYINPUT57), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G1956), .B(n1006), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(KEYINPUT124), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(G1341), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1106 ( .A(KEYINPUT125), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1026), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1029), .Z(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

