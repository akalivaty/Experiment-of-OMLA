//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G169gat), .B(G197gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G229gat), .A2(G233gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G1gat), .B2(new_n211), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(G8gat), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(G50gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(KEYINPUT15), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT88), .B(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n216), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT15), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT14), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT14), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G29gat), .B2(G36gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n225), .B(new_n227), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n219), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n219), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(new_n230), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n233), .A3(new_n234), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n215), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT90), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n231), .B2(new_n215), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  AOI211_X1 g042(.A(KEYINPUT90), .B(new_n215), .C1(new_n236), .C2(new_n238), .ZN(new_n244));
  OAI211_X1 g043(.A(KEYINPUT18), .B(new_n210), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n231), .B(new_n215), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n210), .B(KEYINPUT13), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n239), .A2(new_n240), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n239), .B2(new_n242), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT18), .B1(new_n252), .B2(new_n210), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n209), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n255));
  INV_X1    g054(.A(new_n210), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n238), .ZN(new_n257));
  INV_X1    g056(.A(new_n215), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n241), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n260), .B2(new_n251), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n255), .B1(new_n261), .B2(KEYINPUT18), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n210), .B1(new_n243), .B2(new_n244), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT91), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n249), .A3(new_n208), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n254), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n270));
  OAI21_X1  g069(.A(G120gat), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G120gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G113gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  INV_X1    g075(.A(G127gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n271), .A2(new_n283), .A3(new_n273), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n275), .A2(new_n276), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n290));
  OAI21_X1  g089(.A(G148gat), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n288), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT2), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299));
  INV_X1    g098(.A(G148gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G141gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n295), .A2(new_n298), .B1(new_n288), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT1), .B1(new_n273), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n308));
  OR3_X1    g107(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n285), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT4), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n312));
  INV_X1    g111(.A(new_n273), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT69), .B(G113gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(G120gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n281), .B1(new_n315), .B2(new_n283), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT1), .B1(new_n274), .B2(KEYINPUT70), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n303), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n286), .A2(new_n287), .ZN(new_n321));
  OR2_X1    g120(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n300), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(new_n298), .C1(new_n324), .C2(new_n293), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n302), .A2(new_n288), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n325), .B2(new_n327), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n285), .A2(new_n309), .B1(new_n303), .B2(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n311), .A2(new_n320), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT80), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n311), .A2(new_n320), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n310), .A2(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(new_n332), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n329), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n303), .A2(new_n326), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n318), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n310), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT5), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n337), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G57gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(G85gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n337), .B(new_n352), .C1(new_n341), .C2(new_n347), .ZN(new_n356));
  INV_X1    g155(.A(new_n354), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n339), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n328), .A2(new_n329), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n310), .B1(new_n361), .B2(new_n318), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(new_n335), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n359), .A2(new_n363), .B1(new_n333), .B2(new_n336), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n352), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n355), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  INV_X1    g166(.A(G64gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G92gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT64), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NOR2_X1   g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n379), .A2(new_n381), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n382), .A2(KEYINPUT23), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n386), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT65), .ZN(new_n394));
  AND4_X1   g193(.A1(KEYINPUT25), .A2(new_n392), .A3(new_n385), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n377), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n396), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n376), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n389), .A2(new_n390), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G169gat), .ZN(new_n401));
  INV_X1    g200(.A(G176gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n393), .B1(KEYINPUT26), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT67), .B1(new_n403), .B2(KEYINPUT26), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT67), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n382), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT27), .B(G183gat), .ZN(new_n410));
  INV_X1    g209(.A(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n409), .A2(new_n413), .A3(new_n375), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n373), .B1(new_n400), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G197gat), .B(G204gat), .ZN(new_n419));
  INV_X1    g218(.A(G211gat), .ZN(new_n420));
  INV_X1    g219(.A(G218gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(KEYINPUT22), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G211gat), .B(G218gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n395), .A2(new_n399), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n376), .A2(new_n380), .A3(new_n377), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n380), .B1(new_n376), .B2(new_n377), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n427), .A2(new_n428), .A3(new_n387), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n429), .B2(KEYINPUT25), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n430), .B2(new_n416), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n418), .B(new_n425), .C1(new_n431), .C2(new_n373), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n400), .B2(new_n417), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n372), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n425), .B1(new_n436), .B2(new_n418), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n371), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n418), .B1(new_n431), .B2(new_n373), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n371), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n442), .A4(new_n432), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n433), .A2(new_n437), .A3(new_n371), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n446), .A2(KEYINPUT30), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n438), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n366), .A2(new_n445), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT3), .B1(new_n425), .B2(new_n434), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT82), .B1(new_n451), .B2(new_n303), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n331), .B1(new_n440), .B2(KEYINPUT29), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n325), .A2(new_n327), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n434), .B1(new_n455), .B2(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n440), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n452), .A2(new_n456), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n451), .B2(new_n361), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(G228gat), .A3(G233gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT31), .B(G50gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n466), .A3(new_n462), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n469), .B(G22gat), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n470), .A3(new_n467), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n450), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n352), .B(KEYINPUT83), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n348), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n335), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n310), .C1(new_n361), .C2(new_n318), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT39), .B(new_n481), .C1(new_n333), .C2(new_n480), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n338), .A2(new_n340), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n335), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(new_n477), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n479), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n446), .A2(KEYINPUT30), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n492), .A2(new_n444), .B1(new_n488), .B2(new_n486), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT85), .A2(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(KEYINPUT85), .A2(KEYINPUT38), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n371), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n433), .A2(new_n437), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT37), .B1(new_n441), .B2(new_n432), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n494), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n356), .B(new_n357), .C1(new_n364), .C2(new_n477), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n355), .ZN(new_n502));
  INV_X1    g301(.A(new_n446), .ZN(new_n503));
  INV_X1    g302(.A(new_n496), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n497), .B1(new_n433), .B2(new_n437), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n441), .A2(KEYINPUT37), .A3(new_n432), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n507), .B2(new_n494), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n491), .A2(new_n493), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n476), .B1(new_n509), .B2(new_n475), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n276), .B1(new_n315), .B2(new_n283), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n284), .A2(new_n282), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n309), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n400), .A2(new_n513), .A3(new_n417), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n318), .B1(new_n430), .B2(new_n416), .ZN(new_n515));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(KEYINPUT74), .A3(KEYINPUT34), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n517), .B1(new_n514), .B2(new_n515), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G43gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G71gat), .ZN(new_n526));
  INV_X1    g325(.A(G99gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT33), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(KEYINPUT32), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n524), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT33), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n524), .A2(KEYINPUT71), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n513), .B1(new_n400), .B2(new_n417), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n430), .A2(new_n318), .A3(new_n416), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n516), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n537), .B1(new_n540), .B2(KEYINPUT33), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n524), .A2(KEYINPUT32), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n536), .A2(new_n541), .A3(new_n528), .A4(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n534), .A2(KEYINPUT73), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT73), .B1(new_n534), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n523), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT75), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n534), .A2(new_n522), .A3(new_n543), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(new_n523), .C1(new_n544), .C2(new_n545), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n547), .A2(KEYINPUT36), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n543), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n523), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n548), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n510), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n501), .A2(new_n355), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n492), .A2(new_n444), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n474), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n558), .B1(new_n561), .B2(new_n554), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n547), .A2(new_n548), .A3(new_n550), .A4(new_n474), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n450), .A2(new_n558), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n562), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n268), .B1(new_n557), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT93), .ZN(new_n571));
  INV_X1    g370(.A(G57gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n368), .A2(G57gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT94), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g376(.A(G71gat), .ZN(new_n578));
  INV_X1    g377(.A(G78gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n574), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n576), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n571), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n574), .A2(KEYINPUT95), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n574), .A2(KEYINPUT95), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n573), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n570), .A3(new_n580), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n258), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(G183gat), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n215), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n597));
  INV_X1    g396(.A(G183gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT96), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(G183gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n598), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n600), .A2(G231gat), .A3(G233gat), .A4(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n600), .A2(new_n604), .B1(G231gat), .B2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(new_n420), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n600), .A2(new_n604), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n614), .B2(new_n605), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n593), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n606), .B2(new_n607), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n605), .A3(new_n611), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n592), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n624));
  NAND2_X1  g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT7), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT8), .ZN(new_n627));
  AND2_X1   g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT98), .B(G85gat), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT99), .B(G92gat), .Z(new_n630));
  OAI221_X1 g429(.A(new_n626), .B1(new_n627), .B2(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G99gat), .B(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n628), .A2(new_n627), .ZN(new_n635));
  INV_X1    g434(.A(new_n629), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT99), .B(G92gat), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n632), .A3(new_n626), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n624), .B1(new_n640), .B2(new_n237), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n236), .B2(new_n238), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n642), .A2(G190gat), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n641), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n411), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n421), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(G190gat), .B1(new_n642), .B2(new_n644), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n411), .A3(new_n648), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(G218gat), .A3(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n650), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT101), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n650), .A2(new_n660), .A3(new_n653), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n650), .A2(new_n653), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(new_n656), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT102), .B(new_n657), .C1(new_n650), .C2(new_n653), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n621), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(G230gat), .ZN(new_n669));
  INV_X1    g468(.A(G233gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n589), .A2(new_n639), .A3(new_n634), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n584), .A2(new_n588), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n640), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n643), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(new_n675), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n671), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT103), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G120gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n300), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n676), .A2(new_n677), .ZN(new_n686));
  INV_X1    g485(.A(new_n671), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n679), .A2(new_n671), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n689), .A3(new_n684), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT92), .B(new_n268), .C1(new_n557), .C2(new_n566), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n569), .A2(new_n668), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n366), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n560), .ZN(new_n697));
  NAND2_X1  g496(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n698));
  INV_X1    g497(.A(G8gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n212), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT42), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n699), .B2(new_n697), .ZN(G1325gat));
  INV_X1    g502(.A(G15gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n551), .A2(new_n556), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n694), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n694), .A2(new_n554), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n704), .B2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n694), .A2(new_n474), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  OAI21_X1  g510(.A(new_n667), .B1(new_n557), .B2(new_n566), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT44), .B(new_n667), .C1(new_n557), .C2(new_n566), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n714), .A2(new_n621), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n268), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n691), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n366), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT45), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n569), .A2(new_n621), .A3(new_n692), .A4(new_n693), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n664), .A2(new_n656), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT102), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n664), .A2(new_n663), .A3(new_n656), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(new_n725), .B1(new_n659), .B2(new_n661), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n366), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n223), .A3(new_n728), .ZN(new_n729));
  MUX2_X1   g528(.A(KEYINPUT45), .B(new_n721), .S(new_n729), .Z(G1328gat));
  INV_X1    g529(.A(new_n560), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n224), .A3(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n733));
  OAI21_X1  g532(.A(G36gat), .B1(new_n719), .B2(new_n560), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n705), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n716), .A2(G43gat), .A3(new_n737), .A4(new_n718), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n726), .A3(new_n554), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT104), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n738), .B(new_n742), .C1(new_n739), .C2(G43gat), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT47), .B1(new_n741), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(G1330gat));
  OAI21_X1  g545(.A(new_n220), .B1(new_n719), .B2(new_n474), .ZN(new_n747));
  INV_X1    g546(.A(new_n220), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n748), .A3(new_n475), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g550(.A1(new_n724), .A2(new_n725), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n752), .A2(new_n620), .A3(new_n717), .A4(new_n662), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n692), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT105), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n557), .A2(new_n566), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n728), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n731), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT49), .B(G64gat), .Z(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(G1333gat));
  NOR4_X1   g562(.A1(new_n755), .A2(new_n578), .A3(new_n705), .A4(new_n756), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT106), .ZN(new_n765));
  INV_X1    g564(.A(new_n554), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n757), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n578), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n757), .A2(new_n475), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n714), .A2(new_n715), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n620), .A2(new_n692), .A3(new_n268), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n775), .A2(new_n366), .A3(new_n636), .ZN(new_n776));
  INV_X1    g575(.A(new_n562), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n548), .A2(new_n547), .A3(new_n550), .A4(new_n474), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n564), .ZN(new_n779));
  INV_X1    g578(.A(new_n510), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n705), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n726), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n620), .A2(new_n268), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT51), .A4(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n667), .B(new_n784), .C1(new_n557), .C2(new_n566), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT107), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n785), .A2(new_n788), .B1(new_n787), .B2(new_n786), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n692), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n728), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n776), .B1(new_n791), .B2(new_n636), .ZN(G1336gat));
  INV_X1    g591(.A(new_n786), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n793), .B2(KEYINPUT109), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n794), .A2(new_n796), .B1(new_n788), .B2(new_n785), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n731), .A2(new_n370), .A3(new_n691), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT108), .Z(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n797), .B2(new_n800), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n714), .A2(new_n731), .A3(new_n715), .A4(new_n774), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n630), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n788), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n787), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n801), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT111), .B1(new_n789), .B2(new_n800), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n805), .B(KEYINPUT112), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(new_n817), .B2(new_n630), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n809), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n731), .A4(new_n774), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n630), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n823), .A2(new_n814), .A3(new_n815), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n808), .B1(new_n819), .B2(new_n826), .ZN(G1337gat));
  NOR3_X1   g626(.A1(new_n789), .A2(new_n692), .A3(new_n554), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n737), .A2(G99gat), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(G99gat), .B1(new_n775), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n830), .B(new_n831), .ZN(G1338gat));
  NOR2_X1   g631(.A1(new_n474), .A2(G106gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n798), .A2(new_n691), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G106gat), .B1(new_n775), .B2(new_n474), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n790), .A2(new_n833), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n837), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n836), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(G1339gat));
  NOR2_X1   g639(.A1(new_n753), .A2(new_n691), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n676), .A2(new_n677), .A3(new_n671), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n688), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n684), .B1(new_n678), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n690), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n848), .A2(new_n690), .A3(KEYINPUT115), .A4(new_n849), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n268), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n246), .A2(new_n248), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n243), .A2(new_n244), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n256), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n206), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n691), .C1(new_n267), .C2(new_n266), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n726), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n852), .A2(new_n853), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n267), .B2(new_n266), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n667), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n841), .B1(new_n867), .B2(new_n621), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n731), .A2(new_n366), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n778), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n314), .A3(new_n268), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n868), .B2(new_n475), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n620), .B1(new_n862), .B2(new_n866), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n875), .B(new_n474), .C1(new_n876), .C2(new_n841), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n554), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n870), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n268), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(new_n305), .ZN(G1340gat));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n272), .A3(new_n691), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n691), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(G120gat), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT117), .B(new_n272), .C1(new_n879), .C2(new_n691), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(G1341gat));
  AOI21_X1  g686(.A(G127gat), .B1(new_n872), .B2(new_n620), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n621), .A2(new_n277), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n879), .B2(new_n889), .ZN(G1342gat));
  NOR3_X1   g689(.A1(new_n871), .A2(G134gat), .A3(new_n726), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n879), .A2(new_n667), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n279), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n868), .A2(new_n474), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n737), .A2(new_n366), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT120), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n717), .A2(G141gat), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n901), .A3(new_n897), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n899), .A2(new_n560), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT121), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT119), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n906), .B(new_n907), .C1(new_n868), .C2(new_n474), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n860), .B1(new_n717), .B2(new_n850), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n726), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n620), .B1(new_n910), .B2(new_n866), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT57), .B(new_n475), .C1(new_n911), .C2(new_n841), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n705), .A2(new_n870), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n268), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n289), .A2(new_n290), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR4_X1   g718(.A1(new_n898), .A2(G141gat), .A3(new_n717), .A4(new_n731), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n915), .B2(new_n916), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n904), .A2(new_n919), .B1(new_n918), .B2(new_n921), .ZN(G1344gat));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n726), .A2(new_n850), .A3(new_n864), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n910), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n621), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n726), .A2(new_n620), .A3(new_n692), .A4(new_n717), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT122), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n474), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n924), .B1(new_n930), .B2(KEYINPUT57), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n896), .A2(KEYINPUT57), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n928), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n620), .B1(new_n925), .B2(new_n910), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n475), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(KEYINPUT123), .A3(new_n907), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n691), .A3(new_n914), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n923), .B1(new_n939), .B2(G148gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n913), .A2(new_n691), .A3(new_n914), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(new_n923), .A3(G148gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n899), .A2(new_n560), .A3(new_n902), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n691), .A2(new_n300), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n940), .A2(new_n942), .B1(new_n943), .B2(new_n944), .ZN(G1345gat));
  AND2_X1   g744(.A1(new_n913), .A2(new_n914), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(G155gat), .A3(new_n620), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n296), .B1(new_n943), .B2(new_n621), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1346gat));
  NAND3_X1  g748(.A1(new_n946), .A2(G162gat), .A3(new_n667), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n297), .B1(new_n943), .B2(new_n726), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n728), .A2(new_n560), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n869), .A2(new_n778), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(new_n401), .A3(new_n268), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n953), .B(KEYINPUT124), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n878), .A2(new_n268), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(new_n401), .ZN(G1348gat));
  NAND4_X1  g758(.A1(new_n878), .A2(G176gat), .A3(new_n691), .A4(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n402), .B1(new_n954), .B2(new_n692), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1349gat));
  NAND2_X1  g761(.A1(new_n874), .A2(new_n877), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n963), .A2(new_n620), .A3(new_n766), .A4(new_n957), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n878), .A2(KEYINPUT125), .A3(new_n620), .A4(new_n957), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(G183gat), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n620), .A3(new_n410), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT60), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1350gat));
  NAND3_X1  g773(.A1(new_n955), .A2(new_n411), .A3(new_n667), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n878), .A2(new_n667), .A3(new_n957), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n976), .A2(new_n977), .A3(G190gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n976), .B2(G190gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G1351gat));
  AND2_X1   g779(.A1(new_n705), .A2(new_n957), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n938), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(G197gat), .B1(new_n982), .B2(new_n717), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n896), .A2(new_n705), .A3(new_n953), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n984), .A2(G197gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n717), .B2(new_n985), .ZN(G1352gat));
  NAND3_X1  g785(.A1(new_n938), .A2(new_n691), .A3(new_n981), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G204gat), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n984), .A2(G204gat), .A3(new_n692), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n938), .A2(new_n620), .A3(new_n981), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n620), .A2(new_n420), .ZN(new_n995));
  OAI22_X1  g794(.A1(new_n993), .A2(new_n994), .B1(new_n984), .B2(new_n995), .ZN(G1354gat));
  OAI21_X1  g795(.A(new_n421), .B1(new_n984), .B2(new_n726), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n938), .A2(KEYINPUT127), .A3(new_n981), .ZN(new_n999));
  AND3_X1   g798(.A1(new_n999), .A2(G218gat), .A3(new_n667), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n998), .B1(new_n1000), .B2(new_n1002), .ZN(G1355gat));
endmodule


