//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  XNOR2_X1  g000(.A(KEYINPUT65), .B(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT27), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT27), .B1(new_n206), .B2(KEYINPUT66), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n202), .A2(new_n211), .A3(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT26), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n206), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(new_n214), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n206), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(new_n206), .B2(new_n216), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  AND4_X1   g031(.A1(KEYINPUT25), .A2(new_n230), .A3(new_n218), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n235));
  AOI22_X1  g034(.A1(new_n225), .A2(new_n227), .B1(new_n206), .B2(new_n216), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n218), .A3(new_n232), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT69), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n244), .B(new_n246), .C1(new_n242), .C2(KEYINPUT1), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT68), .B1(new_n248), .B2(new_n249), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n213), .A2(new_n222), .B1(new_n234), .B2(new_n238), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G227gat), .ZN(new_n258));
  INV_X1    g057(.A(G233gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n252), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n250), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n240), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT33), .ZN(new_n265));
  XNOR2_X1  g064(.A(G15gat), .B(G43gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT72), .ZN(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n264), .B(KEYINPUT32), .C1(new_n265), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(KEYINPUT32), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n264), .A2(new_n274), .A3(KEYINPUT32), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n264), .A2(KEYINPUT70), .A3(new_n265), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT70), .B1(new_n264), .B2(new_n265), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n271), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n257), .A2(new_n263), .ZN(new_n281));
  INV_X1    g080(.A(new_n260), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n271), .B(new_n286), .C1(new_n276), .C2(new_n279), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT36), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT36), .B1(new_n288), .B2(new_n289), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G141gat), .B(G148gat), .Z(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n298), .C1(new_n303), .C2(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n311), .B1(G211gat), .B2(G218gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G197gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(G204gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G197gat), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT73), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n313), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G211gat), .B(G218gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n325), .B(new_n313), .C1(new_n316), .C2(new_n321), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(KEYINPUT75), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT75), .B1(new_n324), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n309), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n302), .A2(new_n304), .ZN(new_n331));
  INV_X1    g130(.A(new_n326), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n332), .B2(KEYINPUT85), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n324), .A2(new_n334), .A3(new_n326), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT3), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n330), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G228gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n259), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n326), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n327), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n340), .B1(new_n346), .B2(new_n309), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n324), .B2(new_n326), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n305), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n342), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AND4_X1   g149(.A1(new_n342), .A2(new_n330), .A3(new_n339), .A4(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n341), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G22gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT87), .ZN(new_n354));
  INV_X1    g153(.A(G22gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(new_n341), .C1(new_n350), .C2(new_n351), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G78gat), .B(G106gat), .Z(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT31), .B(G50gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(KEYINPUT87), .A3(G22gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n358), .B(new_n359), .Z(new_n365));
  NAND3_X1  g164(.A1(new_n352), .A2(KEYINPUT88), .A3(G22gat), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n364), .A2(new_n356), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT84), .ZN(new_n370));
  XOR2_X1   g169(.A(G1gat), .B(G29gat), .Z(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G57gat), .B(G85gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n248), .A2(new_n249), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT76), .B1(new_n305), .B2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  AOI211_X1 g180(.A(new_n380), .B(new_n381), .C1(new_n302), .C2(new_n304), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n307), .B(new_n378), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT5), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n262), .A2(new_n388), .A3(new_n389), .A4(new_n331), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n389), .B(new_n331), .C1(new_n251), .C2(new_n252), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n378), .B2(new_n305), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n248), .A2(new_n249), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n331), .A2(new_n395), .A3(KEYINPUT77), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n389), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n387), .B(new_n390), .C1(new_n392), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n331), .A2(new_n395), .A3(KEYINPUT77), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT77), .B1(new_n331), .B2(new_n395), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT4), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n391), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n387), .B1(new_n403), .B2(new_n390), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n386), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n394), .A2(new_n396), .B1(new_n305), .B2(new_n378), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT5), .B1(new_n406), .B2(new_n384), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT79), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n389), .B1(new_n400), .B2(new_n401), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT78), .B1(new_n411), .B2(new_n385), .ZN(new_n412));
  INV_X1    g211(.A(new_n384), .ZN(new_n413));
  INV_X1    g212(.A(new_n379), .ZN(new_n414));
  INV_X1    g213(.A(new_n382), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n306), .A2(new_n395), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n410), .A4(new_n409), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(KEYINPUT5), .C1(new_n406), .C2(new_n384), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n408), .A2(new_n412), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n376), .B(new_n377), .C1(new_n405), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n376), .B1(new_n405), .B2(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(new_n377), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n405), .A2(new_n423), .A3(new_n376), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n240), .A2(new_n308), .B1(G226gat), .B2(G233gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n254), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n346), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n254), .B2(KEYINPUT29), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n240), .A2(G226gat), .A3(G233gat), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n327), .A4(new_n345), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n433), .B2(new_n436), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n433), .A2(new_n436), .ZN(new_n445));
  INV_X1    g244(.A(new_n439), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n370), .B1(new_n429), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n405), .A2(new_n423), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n375), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n428), .A3(new_n377), .ZN(new_n452));
  INV_X1    g251(.A(new_n424), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n448), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n294), .B1(new_n369), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n444), .B2(new_n447), .ZN(new_n460));
  INV_X1    g259(.A(new_n442), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n440), .ZN(new_n462));
  INV_X1    g261(.A(new_n447), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT89), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n425), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n406), .B2(new_n384), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n390), .B1(new_n392), .B2(new_n397), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT82), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n469), .A2(new_n398), .B1(new_n416), .B2(new_n417), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n470), .B2(new_n384), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n383), .B1(new_n399), .B2(new_n404), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n466), .A3(new_n413), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n473), .A3(new_n376), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT40), .A4(new_n376), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n465), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n439), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n445), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n433), .B2(KEYINPUT90), .ZN(new_n484));
  OAI221_X1 g283(.A(new_n479), .B1(new_n442), .B2(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n442), .A2(new_n481), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n433), .B2(new_n436), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT38), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n485), .A2(new_n440), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n452), .A3(new_n453), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n478), .A2(new_n368), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n429), .A2(new_n489), .B1(new_n362), .B2(new_n367), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(KEYINPUT91), .A3(new_n478), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n368), .A2(new_n289), .A3(new_n288), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT35), .B1(new_n457), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n460), .A2(new_n464), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n500), .A2(new_n429), .A3(KEYINPUT35), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(new_n368), .A3(new_n289), .A4(new_n288), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n458), .A2(new_n496), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT12), .ZN(new_n509));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(G1gat), .ZN(new_n512));
  INV_X1    g311(.A(G1gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT16), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n514), .B2(new_n511), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G43gat), .A2(G50gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT94), .B(G43gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(G50gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n522), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT14), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT95), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n521), .A2(new_n523), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n526), .B(new_n528), .C1(new_n524), .C2(new_n525), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT15), .A3(new_n522), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(KEYINPUT96), .A3(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n517), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n533), .A2(KEYINPUT96), .A3(new_n535), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT96), .B1(new_n533), .B2(new_n535), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT17), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n515), .B(G8gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n533), .A2(KEYINPUT17), .A3(new_n535), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n510), .B(new_n540), .C1(new_n543), .C2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n509), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n545), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n517), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n554), .A3(new_n539), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n541), .A2(new_n542), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n553), .A2(new_n555), .B1(new_n556), .B2(new_n517), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n510), .A2(KEYINPUT18), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n544), .B1(new_n541), .B2(new_n542), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n540), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n510), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n551), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n557), .A2(new_n558), .B1(new_n561), .B2(new_n563), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n567), .B(new_n549), .C1(new_n550), .C2(new_n509), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n503), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G57gat), .A2(G64gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(G57gat), .A2(G64gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT100), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G57gat), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577));
  NAND2_X1  g376(.A1(G57gat), .A2(G64gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n579), .A3(KEYINPUT9), .ZN(new_n580));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT9), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT101), .B1(new_n571), .B2(new_n572), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT101), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n576), .A2(new_n589), .A3(new_n578), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G183gat), .B(G211gat), .Z(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  OAI21_X1  g400(.A(new_n544), .B1(new_n593), .B2(new_n592), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT102), .B(KEYINPUT19), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n599), .B(new_n600), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT7), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(G85gat), .ZN(new_n619));
  INV_X1    g418(.A(G92gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(KEYINPUT8), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G99gat), .B(G106gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n617), .B2(new_n621), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n543), .A2(new_n552), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n556), .A2(new_n626), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n610), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n612), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n555), .B(new_n545), .C1(new_n624), .C2(new_n625), .ZN(new_n633));
  INV_X1    g432(.A(new_n612), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n628), .A4(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n632), .A2(new_n639), .A3(new_n635), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n581), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT9), .ZN(new_n645));
  XNOR2_X1  g444(.A(G57gat), .B(G64gat), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(KEYINPUT100), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n647), .B2(new_n579), .ZN(new_n648));
  INV_X1    g447(.A(new_n591), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n648), .A2(new_n649), .B1(new_n624), .B2(new_n625), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n617), .A2(new_n621), .ZN(new_n652));
  INV_X1    g451(.A(new_n622), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n582), .A2(new_n591), .A3(new_n623), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT104), .B1(new_n655), .B2(new_n651), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n646), .A2(KEYINPUT101), .B1(new_n586), .B2(new_n585), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n580), .A2(new_n581), .B1(new_n658), .B2(new_n590), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n626), .A3(new_n660), .A4(KEYINPUT10), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n650), .A2(new_n655), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n667), .A3(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n609), .A2(new_n643), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n454), .A2(KEYINPUT105), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n454), .A2(KEYINPUT105), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n570), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g482(.A1(new_n570), .A2(new_n678), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n516), .B1(new_n685), .B2(new_n500), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n684), .A2(new_n499), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(KEYINPUT42), .B2(new_n688), .ZN(G1325gat));
  OR2_X1    g489(.A1(new_n684), .A2(new_n290), .ZN(new_n691));
  INV_X1    g490(.A(G15gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n294), .B(KEYINPUT106), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT107), .Z(new_n695));
  AOI22_X1  g494(.A1(new_n691), .A2(new_n692), .B1(new_n685), .B2(new_n695), .ZN(G1326gat));
  NOR2_X1   g495(.A1(new_n684), .A2(new_n368), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n503), .B2(new_n643), .ZN(new_n701));
  INV_X1    g500(.A(new_n294), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n429), .A2(new_n370), .A3(new_n448), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT84), .B1(new_n454), .B2(new_n455), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n369), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT91), .B1(new_n494), .B2(new_n478), .ZN(new_n706));
  AND4_X1   g505(.A1(KEYINPUT91), .A2(new_n478), .A3(new_n490), .A4(new_n368), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n702), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n498), .A2(new_n502), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n643), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n609), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n676), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n569), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n681), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n715), .A2(new_n643), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n570), .A2(new_n524), .A3(new_n681), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(G1328gat));
  NAND2_X1  g522(.A1(new_n570), .A2(new_n720), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(G36gat), .A3(new_n499), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n717), .B2(new_n499), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  NAND4_X1  g528(.A1(new_n701), .A2(new_n712), .A3(new_n294), .A4(new_n716), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n520), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n290), .A2(new_n520), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n731), .B(KEYINPUT47), .C1(new_n724), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n724), .A2(new_n732), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n693), .A3(new_n716), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n520), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n724), .B2(new_n368), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n369), .A2(G50gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n717), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n743), .B(new_n739), .C1(new_n717), .C2(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1331gat));
  NAND2_X1  g544(.A1(new_n566), .A2(new_n568), .ZN(new_n746));
  NOR4_X1   g545(.A1(new_n714), .A2(new_n746), .A3(new_n711), .A4(new_n676), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n710), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n681), .A2(KEYINPUT109), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n681), .A2(KEYINPUT109), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n574), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n748), .A2(new_n499), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NOR3_X1   g557(.A1(new_n748), .A2(G71gat), .A3(new_n290), .ZN(new_n759));
  INV_X1    g558(.A(new_n748), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n693), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(G71gat), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1334gat));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n368), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT111), .B(G78gat), .Z(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1335gat));
  NOR3_X1   g566(.A1(new_n609), .A2(new_n746), .A3(new_n676), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n713), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n718), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n609), .A2(new_n746), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n710), .A2(new_n711), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n643), .B1(new_n708), .B2(new_n709), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n681), .A2(new_n619), .A3(new_n675), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n770), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  NOR3_X1   g579(.A1(new_n499), .A2(G92gat), .A3(new_n676), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n701), .A2(new_n712), .A3(new_n500), .A4(new_n768), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n777), .A2(new_n781), .B1(new_n782), .B2(G92gat), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT112), .B1(new_n782), .B2(G92gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n783), .A2(KEYINPUT52), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n776), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n775), .B2(new_n771), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n782), .A2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(KEYINPUT52), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n785), .A2(new_n792), .ZN(G1337gat));
  INV_X1    g592(.A(new_n693), .ZN(new_n794));
  OAI21_X1  g593(.A(G99gat), .B1(new_n769), .B2(new_n794), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n290), .A2(G99gat), .A3(new_n676), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n778), .B2(new_n796), .ZN(G1338gat));
  NOR2_X1   g596(.A1(new_n676), .A2(G106gat), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n369), .B(new_n798), .C1(new_n786), .C2(new_n787), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n701), .A2(new_n712), .A3(new_n369), .A4(new_n768), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n804), .A3(KEYINPUT53), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n799), .B(new_n803), .C1(new_n800), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n678), .A2(new_n569), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n656), .A2(new_n657), .A3(new_n666), .A4(new_n661), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n662), .A2(new_n812), .A3(new_n663), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n672), .A4(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n674), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n813), .A2(new_n672), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n816), .B(KEYINPUT55), .C1(new_n817), .C2(new_n811), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n672), .A3(new_n813), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n815), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n553), .A2(new_n555), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n510), .B1(new_n823), .B2(new_n540), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n561), .A2(new_n563), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n508), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n549), .A2(new_n559), .A3(new_n509), .A4(new_n564), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n641), .A2(new_n642), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n675), .A2(new_n827), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n675), .A2(new_n827), .A3(new_n832), .A4(new_n826), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n831), .B(new_n833), .C1(new_n822), .C2(new_n569), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n829), .B1(new_n834), .B2(new_n643), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n809), .B1(new_n609), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n369), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n718), .A2(new_n500), .A3(new_n290), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n746), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n840), .A2(KEYINPUT116), .A3(G113gat), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT116), .B1(new_n840), .B2(G113gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n751), .A2(new_n837), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n497), .A2(new_n500), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n569), .A2(G113gat), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n841), .A2(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n839), .ZN(new_n848));
  INV_X1    g647(.A(G120gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n676), .ZN(new_n850));
  INV_X1    g649(.A(new_n845), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n675), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n852), .B2(new_n849), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n848), .B2(new_n714), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n714), .A2(G127gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n845), .B2(new_n855), .ZN(G1342gat));
  OR3_X1    g655(.A1(new_n845), .A2(G134gat), .A3(new_n643), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n848), .B2(new_n643), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n749), .A2(new_n750), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT121), .A3(new_n836), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n693), .A2(new_n368), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n864), .A3(new_n499), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT121), .B1(new_n862), .B2(new_n836), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n865), .A2(G141gat), .A3(new_n569), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n702), .A2(new_n499), .A3(new_n681), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n369), .A2(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n677), .A2(new_n746), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n830), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n819), .A2(new_n820), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n746), .A2(new_n815), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n711), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n714), .B1(new_n877), .B2(new_n829), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT118), .B(new_n714), .C1(new_n877), .C2(new_n829), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n871), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n836), .B2(new_n369), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n870), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G141gat), .B1(new_n884), .B2(new_n569), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n876), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n829), .B1(new_n889), .B2(new_n643), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n879), .B1(new_n890), .B2(new_n609), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n881), .A3(new_n809), .ZN(new_n892));
  INV_X1    g691(.A(new_n871), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n822), .A2(new_n569), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n831), .A2(new_n833), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n643), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n829), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n609), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n369), .B1(new_n898), .B2(new_n872), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n892), .A2(new_n893), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT119), .B1(new_n901), .B2(new_n869), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n903), .B(new_n870), .C1(new_n882), .C2(new_n883), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n746), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(G141gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n905), .B2(G141gat), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n907), .A2(new_n908), .A3(new_n867), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n886), .B1(new_n909), .B2(new_n910), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n865), .A2(new_n866), .ZN(new_n912));
  INV_X1    g711(.A(G148gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n675), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n902), .A2(new_n904), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n913), .C1(new_n915), .C2(new_n675), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n872), .B(new_n918), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT57), .B(new_n368), .C1(new_n919), .C2(new_n878), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n900), .B1(new_n836), .B2(new_n369), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n675), .A3(new_n870), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n917), .B1(new_n923), .B2(G148gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n914), .B1(new_n916), .B2(new_n924), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n912), .A2(new_n296), .A3(new_n609), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n915), .A2(new_n609), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n296), .ZN(G1346gat));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n297), .A3(new_n711), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n915), .A2(new_n711), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G162gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1347gat));
  NAND2_X1  g734(.A1(new_n751), .A2(new_n500), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n290), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n838), .ZN(new_n938));
  INV_X1    g737(.A(G169gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(new_n569), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n837), .A2(new_n681), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n497), .A2(new_n499), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G169gat), .B1(new_n944), .B2(new_n746), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n940), .A2(new_n945), .ZN(G1348gat));
  OAI21_X1  g745(.A(G176gat), .B1(new_n938), .B2(new_n676), .ZN(new_n947));
  INV_X1    g746(.A(G176gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n948), .A3(new_n675), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n938), .B2(new_n714), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n941), .A2(new_n211), .A3(new_n943), .A4(new_n609), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n944), .A2(new_n202), .A3(new_n711), .ZN(new_n959));
  OAI21_X1  g758(.A(G190gat), .B1(new_n938), .B2(new_n643), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n936), .A2(new_n693), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n922), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT127), .B1(new_n965), .B2(new_n569), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G197gat), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n965), .A2(KEYINPUT127), .A3(new_n569), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n864), .A2(new_n500), .A3(new_n941), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n746), .A2(new_n317), .ZN(new_n971));
  OAI22_X1  g770(.A1(new_n967), .A2(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1352gat));
  OAI21_X1  g771(.A(G204gat), .B1(new_n965), .B2(new_n676), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n675), .A2(new_n319), .ZN(new_n974));
  OAI21_X1  g773(.A(KEYINPUT62), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  OR3_X1    g774(.A1(new_n969), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n964), .A2(new_n922), .A3(new_n609), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n714), .A2(G211gat), .ZN(new_n981));
  OAI22_X1  g780(.A1(new_n979), .A2(new_n980), .B1(new_n970), .B2(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n965), .B2(new_n643), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n643), .A2(G218gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n970), .B2(new_n984), .ZN(G1355gat));
endmodule


