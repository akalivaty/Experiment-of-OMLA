//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897;
  INV_X1    g000(.A(G1gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G22gat), .Z(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(KEYINPUT16), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(KEYINPUT92), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT93), .B(G8gat), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT93), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(new_n214), .B2(new_n213), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT90), .ZN(new_n217));
  AND2_X1   g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT88), .B(G43gat), .Z(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  AOI211_X1 g019(.A(KEYINPUT15), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT15), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n217), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n213), .B1(new_n228), .B2(new_n212), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n228), .B2(new_n212), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(new_n224), .B2(new_n225), .ZN(new_n231));
  INV_X1    g030(.A(new_n223), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n235));
  AOI21_X1  g034(.A(new_n211), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(KEYINPUT17), .A3(new_n233), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(new_n211), .B2(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n239), .ZN(new_n243));
  INV_X1    g042(.A(new_n211), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(new_n234), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n239), .B(KEYINPUT13), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n242), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n242), .A2(new_n256), .A3(new_n243), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n261));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(KEYINPUT73), .A2(G155gat), .A3(G162gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n267));
  INV_X1    g066(.A(new_n262), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n269));
  INV_X1    g068(.A(G155gat), .ZN(new_n270));
  INV_X1    g069(.A(G162gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n272), .B2(new_n263), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT75), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n262), .B1(new_n276), .B2(KEYINPUT2), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n279));
  INV_X1    g078(.A(G148gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(G141gat), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G148gat), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n277), .A2(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n275), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n280), .A2(KEYINPUT77), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n280), .A2(KEYINPUT77), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n287), .A2(new_n288), .A3(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n280), .B2(G141gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n282), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g092(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n294));
  OAI22_X1  g093(.A1(new_n289), .A2(new_n293), .B1(new_n268), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n285), .A2(new_n286), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT22), .ZN(new_n300));
  INV_X1    g099(.A(G211gat), .ZN(new_n301));
  INV_X1    g100(.A(G218gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G211gat), .B(G218gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n284), .B1(new_n274), .B2(new_n273), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n295), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n286), .B1(new_n306), .B2(KEYINPUT29), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n298), .A2(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT84), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT31), .B(G50gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(G22gat), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n311), .B(new_n312), .Z(new_n320));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G22gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n323), .B(new_n317), .C1(new_n313), .C2(KEYINPUT84), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n319), .B2(new_n324), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n261), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n327), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT85), .A3(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  INV_X1    g135(.A(G120gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G113gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  INV_X1    g139(.A(G134gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G127gat), .ZN(new_n342));
  INV_X1    g141(.A(G127gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G134gat), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n339), .A2(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n344), .A3(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(KEYINPUT66), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G120gat), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n347), .A2(new_n349), .A3(G113gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n350), .B2(KEYINPUT67), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT66), .B(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n336), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n345), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n309), .B2(KEYINPUT3), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT5), .B(new_n334), .C1(new_n357), .C2(new_n296), .ZN(new_n358));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n268), .B1(new_n278), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n291), .A2(new_n292), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT77), .B(G148gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G141gat), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G141gat), .B(G148gat), .Z(new_n365));
  NAND2_X1  g164(.A1(new_n276), .A2(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n278), .A2(KEYINPUT75), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n262), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n266), .A2(KEYINPUT74), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n364), .B1(new_n369), .B2(new_n275), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .A4(new_n356), .ZN(new_n373));
  INV_X1    g172(.A(new_n345), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n352), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n346), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n336), .A2(new_n354), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n350), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n374), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT4), .B1(new_n309), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n356), .A2(new_n372), .A3(new_n295), .A4(new_n285), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(KEYINPUT79), .A3(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n358), .A2(KEYINPUT80), .A3(new_n373), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n373), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n370), .B2(new_n286), .ZN(new_n388));
  INV_X1    g187(.A(new_n296), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n387), .B(new_n333), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n385), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n382), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n357), .A2(new_n296), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(KEYINPUT4), .C1(new_n309), .C2(new_n380), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n333), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n309), .A2(new_n380), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n356), .A2(new_n295), .A3(new_n285), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n387), .B1(new_n404), .B2(new_n334), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT6), .B1(new_n392), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408));
  INV_X1    g207(.A(new_n396), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n384), .A2(new_n391), .B1(new_n401), .B2(new_n405), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT81), .B(KEYINPUT6), .C1(new_n392), .C2(new_n406), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT82), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n333), .B(new_n400), .C1(new_n388), .C2(new_n389), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n382), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n409), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n391), .B2(new_n384), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT81), .B1(new_n418), .B2(KEYINPUT6), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n407), .A2(new_n408), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n410), .A2(new_n409), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n413), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT27), .B(G183gat), .ZN(new_n427));
  INV_X1    g226(.A(G190gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT28), .ZN(new_n430));
  NAND2_X1  g229(.A1(G169gat), .A2(G176gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT26), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n435));
  INV_X1    g234(.A(G183gat), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n434), .A2(new_n435), .B1(new_n436), .B2(new_n428), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n432), .A2(KEYINPUT23), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT65), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n436), .A2(new_n428), .A3(KEYINPUT24), .ZN(new_n441));
  XOR2_X1   g240(.A(G183gat), .B(G190gat), .Z(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT24), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT64), .B(G169gat), .ZN(new_n444));
  INV_X1    g243(.A(G176gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT23), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n440), .A2(new_n443), .A3(new_n431), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n431), .A2(KEYINPUT25), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(KEYINPUT23), .B2(new_n432), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n440), .A2(new_n443), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n438), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n453), .B2(KEYINPUT29), .ZN(new_n456));
  INV_X1    g255(.A(new_n306), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n455), .B2(new_n456), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G8gat), .B(G36gat), .Z(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT71), .ZN(new_n463));
  XOR2_X1   g262(.A(G64gat), .B(G92gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(KEYINPUT72), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n460), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n466), .A3(new_n458), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT72), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n467), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT70), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(KEYINPUT70), .A3(new_n458), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI22_X1  g276(.A1(new_n477), .A2(new_n466), .B1(new_n472), .B2(new_n469), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n426), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT83), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n426), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n332), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n453), .B(new_n380), .ZN(new_n486));
  NAND2_X1  g285(.A1(G227gat), .A2(G233gat), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT32), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT69), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT32), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G43gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(G71gat), .B(G99gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n488), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n487), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n499), .B(KEYINPUT34), .Z(new_n500));
  OAI211_X1 g299(.A(new_n488), .B(KEYINPUT32), .C1(new_n496), .C2(new_n495), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n500), .B1(new_n498), .B2(new_n501), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n485), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(KEYINPUT36), .A3(new_n502), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n260), .B1(new_n484), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n483), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n482), .B1(new_n426), .B2(new_n479), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n331), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT86), .A3(new_n508), .ZN(new_n514));
  INV_X1    g313(.A(new_n479), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n383), .A2(new_n373), .A3(new_n398), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n334), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(KEYINPUT39), .C1(new_n334), .C2(new_n404), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(new_n409), .C1(KEYINPUT39), .C2(new_n517), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT40), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n422), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n329), .A2(new_n325), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n422), .A2(new_n424), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n407), .B2(new_n422), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n467), .A2(new_n471), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT37), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n466), .B1(new_n461), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n477), .B2(new_n528), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT38), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT38), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n529), .B(new_n532), .C1(new_n528), .C2(new_n461), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n525), .A2(new_n527), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n521), .A2(new_n523), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n510), .A2(new_n514), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n506), .A2(new_n502), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n481), .A2(new_n538), .A3(new_n483), .A4(new_n523), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n479), .A2(new_n541), .ZN(new_n542));
  NOR4_X1   g341(.A1(new_n537), .A2(new_n542), .A3(new_n522), .A4(new_n525), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n259), .B1(new_n536), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  XOR2_X1   g347(.A(G57gat), .B(G64gat), .Z(new_n549));
  AOI211_X1 g348(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(KEYINPUT9), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(KEYINPUT9), .B2(new_n548), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT94), .B(G57gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G64gat), .ZN(new_n553));
  INV_X1    g352(.A(G64gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G57gat), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G127gat), .B(G155gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT95), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G183gat), .B(G211gat), .Z(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  OAI21_X1  g365(.A(new_n244), .B1(new_n558), .B2(new_n557), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n566), .B(new_n569), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n234), .A2(new_n235), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT7), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n579), .B(KEYINPUT97), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n237), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n234), .A2(new_n589), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT96), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n571), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n587), .A2(new_n557), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT98), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n557), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n587), .A2(KEYINPUT98), .A3(new_n557), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT10), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n605), .A2(KEYINPUT10), .ZN(new_n611));
  INV_X1    g410(.A(G230gat), .ZN(new_n612));
  INV_X1    g411(.A(G233gat), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(new_n615), .A3(new_n609), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n614), .B2(new_n616), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n604), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n426), .A2(KEYINPUT99), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n426), .A2(KEYINPUT99), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n546), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g430(.A1(new_n546), .A2(new_n625), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n479), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n634), .A2(KEYINPUT100), .B1(KEYINPUT42), .B2(new_n209), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(KEYINPUT100), .B2(new_n634), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT16), .B(G8gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n641), .ZN(G1325gat));
  OAI21_X1  g441(.A(G15gat), .B1(new_n632), .B2(new_n508), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n537), .A2(G15gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n632), .B2(new_n644), .ZN(G1326gat));
  NAND3_X1  g444(.A1(new_n546), .A2(new_n331), .A3(new_n625), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT102), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT43), .B(G22gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  AND4_X1   g448(.A1(new_n546), .A2(new_n570), .A3(new_n602), .A4(new_n623), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n224), .A3(new_n629), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT45), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n513), .A2(new_n508), .A3(new_n535), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n545), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n602), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n603), .B1(new_n536), .B2(new_n545), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n659), .A2(new_n258), .A3(new_n570), .A4(new_n623), .ZN(new_n660));
  OAI21_X1  g459(.A(G29gat), .B1(new_n660), .B2(new_n628), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n661), .ZN(G1328gat));
  NAND3_X1  g461(.A1(new_n650), .A2(new_n225), .A3(new_n515), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT46), .Z(new_n664));
  OAI21_X1  g463(.A(G36gat), .B1(new_n660), .B2(new_n479), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(new_n660), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n219), .B1(new_n667), .B2(new_n509), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n538), .A2(new_n219), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n650), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g470(.A1(new_n650), .A2(new_n220), .A3(new_n331), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT48), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n522), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(G50gat), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  OAI21_X1  g477(.A(G50gat), .B1(new_n660), .B2(new_n332), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n679), .A2(new_n672), .ZN(new_n680));
  OAI22_X1  g479(.A1(new_n677), .A2(new_n678), .B1(KEYINPUT48), .B2(new_n680), .ZN(G1331gat));
  NOR3_X1   g480(.A1(new_n604), .A2(new_n258), .A3(new_n623), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n654), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n629), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(new_n552), .Z(G1332gat));
  INV_X1    g484(.A(KEYINPUT49), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n515), .B1(new_n686), .B2(new_n554), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT105), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n554), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1333gat));
  NAND2_X1  g490(.A1(new_n683), .A2(new_n509), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n537), .A2(G71gat), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n692), .A2(G71gat), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1334gat));
  NAND2_X1  g495(.A1(new_n683), .A2(new_n331), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT107), .B(G78gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1335gat));
  NOR2_X1   g498(.A1(new_n571), .A2(new_n258), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n623), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n659), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n659), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G85gat), .B1(new_n707), .B2(new_n628), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n603), .B1(new_n545), .B2(new_n653), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n701), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n711), .B(KEYINPUT51), .C1(new_n710), .C2(new_n709), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  INV_X1    g512(.A(new_n653), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n543), .B1(new_n539), .B2(KEYINPUT35), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n602), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n700), .B1(new_n716), .B2(KEYINPUT109), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n709), .A2(new_n710), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT110), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(KEYINPUT110), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n624), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n629), .A2(new_n576), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n708), .B1(new_n723), .B2(new_n724), .ZN(G1336gat));
  OAI21_X1  g524(.A(G92gat), .B1(new_n703), .B2(new_n479), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n623), .A2(G92gat), .A3(new_n479), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT111), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n726), .B(new_n727), .C1(new_n720), .C2(new_n729), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n659), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT108), .B1(new_n659), .B2(new_n702), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n731), .A2(new_n732), .A3(new_n479), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n733), .A2(new_n577), .B1(new_n720), .B2(new_n729), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT112), .B1(new_n734), .B2(KEYINPUT52), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n729), .B1(new_n712), .B2(new_n719), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n705), .A2(new_n515), .A3(new_n706), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n738), .A2(new_n739), .A3(new_n727), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n730), .B1(new_n735), .B2(new_n740), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n707), .B2(new_n508), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n537), .A2(G99gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n723), .B2(new_n743), .ZN(G1338gat));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT113), .B(G106gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n703), .B2(new_n523), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n623), .A2(new_n523), .A3(G106gat), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n745), .B(new_n747), .C1(new_n720), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n720), .A2(new_n748), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n705), .A2(new_n331), .A3(new_n706), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n746), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n752), .B2(new_n745), .ZN(G1339gat));
  NAND2_X1  g552(.A1(new_n625), .A2(new_n259), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n610), .A2(new_n611), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n615), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(KEYINPUT54), .A3(new_n614), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n614), .A2(KEYINPUT54), .ZN(new_n758));
  INV_X1    g557(.A(new_n619), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT55), .A4(new_n759), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n620), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT114), .B1(new_n238), .B2(new_n239), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n245), .A2(new_n247), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n238), .A2(KEYINPUT114), .A3(new_n239), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n253), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n257), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n764), .A2(new_n603), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n762), .A2(new_n258), .A3(new_n620), .A4(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n623), .B2(new_n770), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n603), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n754), .B1(new_n774), .B2(new_n571), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(new_n538), .A3(new_n332), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n628), .A2(new_n515), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G113gat), .B1(new_n778), .B2(new_n259), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n775), .A2(new_n629), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n780), .A2(new_n479), .A3(new_n538), .A4(new_n523), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT115), .Z(new_n782));
  NAND2_X1  g581(.A1(new_n258), .A2(new_n335), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(G1340gat));
  NAND2_X1  g583(.A1(new_n624), .A2(new_n352), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n776), .A2(new_n624), .A3(new_n777), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n786), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT116), .B1(new_n786), .B2(G120gat), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n782), .A2(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G1341gat));
  OAI21_X1  g588(.A(G127gat), .B1(new_n778), .B2(new_n570), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n571), .A2(new_n343), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT117), .Z(G1342gat));
  NOR3_X1   g592(.A1(new_n603), .A2(G134gat), .A3(new_n515), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n780), .A2(new_n538), .A3(new_n523), .A4(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n795), .A2(KEYINPUT56), .ZN(new_n796));
  OAI21_X1  g595(.A(G134gat), .B1(new_n778), .B2(new_n603), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(KEYINPUT56), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT118), .Z(G1343gat));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n522), .A3(new_n508), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n515), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n259), .A2(G141gat), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT58), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n623), .A2(new_n770), .A3(KEYINPUT120), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT120), .B1(new_n623), .B2(new_n770), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n772), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n602), .B1(new_n808), .B2(new_n809), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n771), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n754), .B1(new_n812), .B2(new_n571), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n805), .B1(new_n813), .B2(new_n331), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n777), .A2(new_n508), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT119), .Z(new_n816));
  NAND2_X1  g615(.A1(new_n775), .A2(new_n522), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(KEYINPUT57), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n259), .ZN(new_n820));
  OAI21_X1  g619(.A(G141gat), .B1(new_n820), .B2(KEYINPUT122), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT122), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n819), .A2(new_n822), .A3(new_n259), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n804), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n802), .A2(new_n803), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n820), .B2(new_n282), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT58), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(G1344gat));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n819), .A2(new_n623), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n362), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n802), .A2(new_n362), .A3(new_n624), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n813), .B2(new_n331), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n833), .A2(new_n834), .B1(new_n817), .B2(new_n805), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n816), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n623), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n831), .B(new_n832), .C1(new_n839), .C2(new_n840), .ZN(G1345gat));
  OAI21_X1  g640(.A(G155gat), .B1(new_n819), .B2(new_n570), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n802), .A2(new_n270), .A3(new_n571), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1346gat));
  OAI21_X1  g643(.A(G162gat), .B1(new_n819), .B2(new_n603), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n602), .A2(new_n271), .A3(new_n479), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n801), .B2(new_n846), .ZN(G1347gat));
  AND2_X1   g646(.A1(new_n775), .A2(new_n628), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n515), .A2(new_n848), .A3(new_n538), .A4(new_n523), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n258), .A3(new_n444), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n629), .A2(new_n479), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n776), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G169gat), .B1(new_n852), .B2(new_n259), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT124), .ZN(G1348gat));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n445), .A3(new_n624), .ZN(new_n856));
  OAI21_X1  g655(.A(G176gat), .B1(new_n852), .B2(new_n623), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1349gat));
  AND2_X1   g657(.A1(new_n571), .A2(new_n427), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n849), .A2(new_n859), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n860));
  OAI21_X1  g659(.A(G183gat), .B1(new_n852), .B2(new_n570), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n862), .B(new_n863), .Z(G1350gat));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n428), .A3(new_n602), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n776), .A2(new_n602), .A3(new_n851), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n868));
  AND4_X1   g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(G190gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n428), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n867), .A2(new_n870), .B1(new_n866), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n869), .B2(new_n871), .ZN(G1351gat));
  NOR3_X1   g671(.A1(new_n509), .A2(new_n479), .A3(new_n523), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(G197gat), .B1(new_n875), .B2(new_n258), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n835), .A2(new_n836), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n629), .A2(new_n509), .A3(new_n479), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n258), .A2(G197gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(G1352gat));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n624), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G204gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n874), .A2(G204gat), .A3(new_n623), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(KEYINPUT127), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n883), .A2(new_n886), .A3(new_n888), .ZN(G1353gat));
  NAND3_X1  g688(.A1(new_n875), .A2(new_n301), .A3(new_n571), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n571), .B(new_n878), .C1(new_n835), .C2(new_n836), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT63), .B1(new_n891), .B2(G211gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1354gat));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n302), .A3(new_n602), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n602), .A3(new_n878), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n302), .ZN(G1355gat));
endmodule


