//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G227gat), .ZN(new_n205));
  INV_X1    g004(.A(G233gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G113gat), .B2(G120gat), .ZN(new_n221));
  AND2_X1   g020(.A1(G113gat), .A2(G120gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n216), .A2(new_n219), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n211), .B(new_n224), .C1(new_n230), .C2(new_n209), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n215), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n222), .B2(new_n221), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n227), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT24), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(G183gat), .ZN(new_n243));
  INV_X1    g042(.A(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(G169gat), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT25), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n250), .A2(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n246), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(KEYINPUT23), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n250), .B1(G169gat), .B2(G176gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n258), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n261), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n237), .A2(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT25), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT26), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n257), .A2(new_n258), .B1(new_n269), .B2(new_n253), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n236), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n243), .A2(KEYINPUT27), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT27), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G183gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n280), .A3(new_n244), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n277), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n244), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n276), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n235), .A2(new_n268), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n267), .A3(new_n260), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n231), .A2(new_n227), .A3(new_n233), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n208), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n204), .B1(new_n295), .B2(KEYINPUT33), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n289), .A2(new_n294), .ZN(new_n300));
  AOI221_X4 g099(.A(new_n297), .B1(KEYINPUT33), .B2(new_n204), .C1(new_n300), .C2(new_n207), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n290), .A2(new_n293), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n290), .A2(new_n293), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT73), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n307), .A3(new_n294), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n308), .A3(new_n208), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n300), .A2(KEYINPUT34), .A3(new_n207), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n303), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n309), .A2(new_n314), .A3(new_n311), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n309), .B2(new_n311), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n303), .B(new_n317), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n302), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G22gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G228gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(KEYINPUT81), .A3(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(G141gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G148gat), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G141gat), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n335), .A2(new_n337), .B1(KEYINPUT2), .B2(new_n329), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n331), .B(new_n330), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G211gat), .ZN(new_n345));
  INV_X1    g144(.A(G218gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G211gat), .A2(G218gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G197gat), .B(G204gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT22), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(KEYINPUT76), .A3(new_n348), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G211gat), .B(G218gat), .Z(new_n358));
  NOR3_X1   g157(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT77), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n360));
  INV_X1    g159(.A(G197gat), .ZN(new_n361));
  INV_X1    g160(.A(G204gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n363), .A2(new_n364), .B1(new_n353), .B2(new_n348), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n360), .B1(new_n365), .B2(new_n349), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n357), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n344), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n367), .B(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n343), .A2(new_n371), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n369), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n325), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n367), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n325), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT77), .B1(new_n355), .B2(new_n358), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n365), .A2(new_n360), .A3(new_n349), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n383), .A2(new_n384), .B1(new_n358), .B2(new_n355), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n369), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT84), .B1(new_n385), .B2(KEYINPUT29), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n371), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n382), .B1(new_n344), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n324), .B1(new_n379), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT86), .ZN(new_n393));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n344), .ZN(new_n397));
  INV_X1    g196(.A(new_n382), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n373), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n371), .A3(new_n370), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n401), .A2(new_n344), .B1(new_n375), .B2(new_n377), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n399), .B(G22gat), .C1(new_n402), .C2(new_n325), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n393), .A2(new_n396), .B1(new_n392), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405));
  AND4_X1   g204(.A1(new_n405), .A2(new_n403), .A3(new_n392), .A4(new_n396), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n207), .B1(new_n304), .B2(new_n305), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(new_n204), .C1(KEYINPUT33), .C2(new_n295), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n296), .A2(new_n298), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT71), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT71), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n416), .A3(new_n321), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n290), .B2(new_n369), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n268), .B2(new_n288), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n375), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n290), .A2(new_n369), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n422), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n290), .A2(new_n423), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n367), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n424), .A2(new_n425), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n433), .B2(new_n367), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n421), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT80), .B(new_n421), .C1(new_n432), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n339), .A2(KEYINPUT3), .A3(new_n342), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n376), .A2(new_n225), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n343), .A2(new_n233), .A3(new_n231), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n235), .A2(new_n343), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n447), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n447), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n291), .A2(new_n343), .A3(KEYINPUT4), .A4(new_n292), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n441), .A2(new_n452), .A3(new_n442), .A4(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n225), .A2(new_n339), .A3(new_n342), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n442), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n443), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT0), .ZN(new_n462));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n460), .A2(new_n465), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n445), .A2(new_n450), .B1(new_n454), .B2(new_n458), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n466), .B1(new_n470), .B2(new_n464), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n468), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n428), .A2(new_n430), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT79), .B1(new_n473), .B2(new_n380), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(new_n426), .A3(new_n431), .A4(new_n420), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT30), .ZN(new_n476));
  INV_X1    g275(.A(new_n432), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n474), .A4(new_n420), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n439), .A2(new_n472), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n323), .A2(new_n407), .A3(new_n417), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n486));
  INV_X1    g285(.A(new_n302), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n416), .A2(new_n487), .A3(new_n321), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n323), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n393), .A2(new_n396), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n403), .A2(new_n392), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n403), .A2(new_n392), .A3(new_n405), .A4(new_n396), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n437), .A2(new_n438), .B1(new_n476), .B2(new_n479), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n472), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n323), .A2(KEYINPUT89), .A3(new_n488), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n491), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n414), .A2(new_n416), .A3(new_n321), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n487), .B1(new_n416), .B2(new_n321), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT36), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n323), .A2(new_n507), .A3(new_n488), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n435), .B1(new_n510), .B2(new_n420), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n477), .B2(new_n474), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT38), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n468), .B(new_n475), .C1(new_n469), .C2(new_n471), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n473), .A2(KEYINPUT88), .A3(new_n375), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT88), .B1(new_n473), .B2(new_n375), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n516), .B(new_n517), .C1(new_n367), .C2(new_n433), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT38), .B1(new_n518), .B2(KEYINPUT37), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n511), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n496), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT40), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n450), .A2(new_n441), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n457), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n464), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n446), .A2(new_n442), .A3(new_n455), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT39), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n523), .B2(new_n457), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n522), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(KEYINPUT40), .A3(new_n464), .A4(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n460), .A2(new_n465), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(new_n497), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT87), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n534), .A2(new_n497), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n521), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n496), .A2(new_n498), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n509), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n503), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT93), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G1gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n544), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n545), .A3(G1gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G29gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n564));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(KEYINPUT17), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n566), .B2(new_n567), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n555), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n554), .A3(new_n568), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n576));
  INV_X1    g375(.A(new_n568), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n574), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n573), .B(KEYINPUT13), .Z(new_n580));
  AOI22_X1  g379(.A1(new_n575), .A2(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n572), .A2(KEYINPUT18), .A3(new_n573), .A4(new_n574), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT12), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n581), .A2(new_n582), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(KEYINPUT95), .A3(new_n592), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n542), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT97), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n326), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G57gat), .A2(G64gat), .ZN(new_n604));
  OR2_X1    g403(.A1(G57gat), .A2(G64gat), .ZN(new_n605));
  INV_X1    g404(.A(G71gat), .ZN(new_n606));
  INV_X1    g405(.A(G78gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n604), .B(new_n605), .C1(new_n608), .C2(KEYINPUT9), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT96), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n607), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n612), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(new_n214), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n553), .A2(new_n554), .B1(KEYINPUT21), .B2(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(G127gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n603), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n625), .A3(new_n603), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT100), .ZN(new_n631));
  OR2_X1    g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633));
  NAND2_X1  g432(.A1(G99gat), .A2(G106gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT8), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n634), .B2(KEYINPUT99), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(KEYINPUT99), .B2(new_n634), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT7), .ZN(new_n640));
  INV_X1    g439(.A(G85gat), .ZN(new_n641));
  OAI21_X1  g440(.A(G92gat), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n642), .A2(new_n644), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n636), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n639), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n635), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n568), .A2(new_n650), .B1(KEYINPUT41), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n569), .A2(new_n571), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n650), .ZN(new_n655));
  XOR2_X1   g454(.A(G190gat), .B(G218gat), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT98), .Z(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n656), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n653), .B(new_n664), .C1(new_n654), .C2(new_n650), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n657), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n661), .B(new_n662), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n657), .B2(new_n665), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n636), .A2(KEYINPUT102), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n615), .A2(new_n646), .A3(new_n649), .A4(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n613), .A3(new_n614), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT10), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n650), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n676));
  INV_X1    g475(.A(G230gat), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n675), .A2(new_n676), .B1(new_n677), .B2(new_n206), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n206), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n678), .A2(new_n680), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n629), .A2(new_n670), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n598), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n472), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  INV_X1    g493(.A(new_n497), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G8gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n548), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n691), .B2(new_n695), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT42), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT42), .B2(new_n700), .ZN(G1325gat));
  INV_X1    g502(.A(new_n691), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n704), .B2(new_n509), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n491), .A2(new_n501), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n704), .B2(new_n707), .ZN(G1326gat));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n496), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT43), .B(G22gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  INV_X1    g512(.A(new_n597), .ZN(new_n714));
  INV_X1    g513(.A(new_n629), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n669), .A3(new_n689), .ZN(new_n716));
  AOI211_X1 g515(.A(new_n714), .B(new_n716), .C1(new_n503), .C2(new_n541), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n692), .A2(new_n560), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n713), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n716), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n542), .A2(new_n597), .A3(new_n721), .A4(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(KEYINPUT103), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n712), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n717), .A2(new_n713), .A3(new_n719), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(KEYINPUT103), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n627), .A2(KEYINPUT104), .A3(new_n628), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n730));
  INV_X1    g529(.A(new_n628), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n626), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n581), .A2(new_n582), .A3(new_n589), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n589), .B1(new_n581), .B2(new_n582), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n733), .A2(new_n736), .A3(new_n688), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n542), .A2(KEYINPUT105), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n503), .A2(new_n541), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n670), .A2(KEYINPUT44), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n542), .A2(new_n669), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n738), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n560), .B1(new_n746), .B2(new_n692), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT106), .B1(new_n728), .B2(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n503), .A2(new_n740), .A3(new_n541), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n740), .B1(new_n503), .B2(new_n541), .ZN(new_n750));
  INV_X1    g549(.A(new_n742), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n542), .B2(new_n669), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n692), .B(new_n737), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G29gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n756), .A2(new_n757), .A3(new_n727), .A4(new_n724), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n748), .A2(new_n758), .ZN(G1328gat));
  NAND3_X1  g558(.A1(new_n717), .A2(new_n556), .A3(new_n695), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT46), .Z(new_n761));
  AND2_X1   g560(.A1(new_n746), .A2(new_n695), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n556), .ZN(G1329gat));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764));
  INV_X1    g563(.A(G43gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n506), .A2(new_n508), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n746), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n717), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n768), .A2(G43gat), .A3(new_n706), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n769), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n509), .B(new_n738), .C1(new_n743), .C2(new_n745), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT47), .B(new_n771), .C1(new_n772), .C2(new_n765), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1330gat));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n746), .B2(new_n496), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n768), .A2(G50gat), .A3(new_n407), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n778), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n407), .B(new_n738), .C1(new_n743), .C2(new_n745), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT48), .B(new_n780), .C1(new_n781), .C2(new_n776), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1331gat));
  NOR2_X1   g582(.A1(new_n749), .A2(new_n750), .ZN(new_n784));
  NOR4_X1   g583(.A1(new_n715), .A2(new_n593), .A3(new_n669), .A4(new_n689), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n692), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g588(.A(new_n497), .B(KEYINPUT107), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT49), .B(G64gat), .Z(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(G1333gat));
  OAI21_X1  g594(.A(G71gat), .B1(new_n786), .B2(new_n509), .ZN(new_n796));
  INV_X1    g595(.A(new_n706), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n606), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n786), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n796), .B(KEYINPUT50), .C1(new_n786), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1334gat));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n407), .ZN(new_n804));
  XNOR2_X1  g603(.A(KEYINPUT108), .B(G78gat), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1335gat));
  NOR2_X1   g605(.A1(new_n629), .A2(new_n593), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n542), .A2(new_n669), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT51), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n811), .A2(KEYINPUT109), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(KEYINPUT109), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n641), .A3(new_n692), .A4(new_n688), .ZN(new_n816));
  INV_X1    g615(.A(new_n807), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n689), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n752), .B2(new_n754), .ZN(new_n819));
  OAI21_X1  g618(.A(G85gat), .B1(new_n819), .B2(new_n472), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(G1336gat));
  NAND3_X1  g620(.A1(new_n791), .A2(new_n643), .A3(new_n688), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT110), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n810), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  INV_X1    g624(.A(new_n818), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n790), .B(new_n826), .C1(new_n743), .C2(new_n745), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n824), .B(new_n825), .C1(new_n827), .C2(new_n643), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n808), .A2(new_n829), .A3(KEYINPUT51), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT51), .B1(new_n808), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n695), .B(new_n818), .C1(new_n752), .C2(new_n754), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n823), .A2(new_n832), .B1(new_n833), .B2(G92gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n828), .B1(new_n834), .B2(new_n825), .ZN(G1337gat));
  NOR3_X1   g634(.A1(new_n706), .A2(G99gat), .A3(new_n689), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n815), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G99gat), .B1(new_n819), .B2(new_n509), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1338gat));
  OAI211_X1 g638(.A(new_n496), .B(new_n818), .C1(new_n752), .C2(new_n754), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G106gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n407), .A2(G106gat), .A3(new_n689), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n810), .A2(new_n814), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n832), .A2(new_n843), .B1(new_n840), .B2(G106gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n842), .ZN(G1339gat));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n848));
  INV_X1    g647(.A(new_n580), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n578), .A2(new_n574), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT112), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n578), .A2(new_n852), .A3(new_n574), .A4(new_n849), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n572), .A2(new_n574), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n851), .B(new_n853), .C1(new_n854), .C2(new_n573), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n588), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n592), .A3(new_n688), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n675), .A2(new_n676), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n679), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n860), .A2(KEYINPUT54), .A3(new_n678), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n685), .B1(new_n678), .B2(KEYINPUT54), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(KEYINPUT54), .A3(new_n678), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n678), .A2(KEYINPUT54), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT55), .A4(new_n685), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n687), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n857), .B1(new_n867), .B2(new_n736), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n670), .ZN(new_n869));
  INV_X1    g668(.A(new_n867), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT113), .B1(new_n856), .B2(new_n592), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n856), .A2(KEYINPUT113), .A3(new_n592), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n870), .A2(new_n872), .A3(new_n669), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n733), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n690), .A2(new_n593), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n848), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n729), .A2(new_n732), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n593), .A2(new_n687), .A3(new_n866), .A4(new_n863), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n669), .B1(new_n879), .B2(new_n857), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n669), .A2(new_n863), .A3(new_n687), .A4(new_n866), .ZN(new_n881));
  INV_X1    g680(.A(new_n873), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n881), .A2(new_n882), .A3(new_n871), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n690), .A2(new_n593), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(KEYINPUT114), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n504), .A2(new_n496), .A3(new_n505), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n877), .A2(new_n886), .A3(new_n692), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n791), .ZN(new_n889));
  AOI21_X1  g688(.A(G113gat), .B1(new_n889), .B2(new_n593), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n797), .A2(new_n692), .A3(new_n790), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n877), .A2(new_n886), .A3(new_n407), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n886), .A3(KEYINPUT115), .A4(new_n407), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n714), .A2(new_n209), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(G1340gat));
  NAND3_X1  g697(.A1(new_n889), .A2(new_n230), .A3(new_n688), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n688), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT116), .B1(new_n900), .B2(G120gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1341gat));
  NAND3_X1  g702(.A1(new_n889), .A2(new_n214), .A3(new_n629), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n896), .A2(new_n733), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n214), .ZN(G1342gat));
  AOI21_X1  g705(.A(new_n212), .B1(new_n896), .B2(new_n669), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n695), .A2(new_n670), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n212), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n888), .A2(KEYINPUT56), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT56), .B1(new_n888), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n907), .A2(KEYINPUT117), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT117), .B1(new_n907), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1343gat));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n857), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n856), .A2(KEYINPUT118), .A3(new_n592), .A4(new_n688), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n866), .A2(new_n687), .ZN(new_n920));
  INV_X1    g719(.A(new_n862), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n864), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT55), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(KEYINPUT119), .A3(new_n864), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n919), .B1(new_n597), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n874), .B1(new_n927), .B2(new_n669), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n876), .B1(new_n928), .B2(new_n715), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT57), .B1(new_n929), .B2(new_n407), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n877), .A2(new_n886), .A3(new_n931), .A4(new_n496), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n766), .A2(new_n472), .A3(new_n791), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G141gat), .B1(new_n934), .B2(new_n714), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n877), .A2(new_n886), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n766), .A2(new_n407), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n692), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n791), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n597), .A2(new_n334), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT120), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT58), .B1(new_n935), .B2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT58), .B(G141gat), .C1(new_n934), .C2(new_n736), .ZN(new_n945));
  NOR2_X1   g744(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n939), .B2(new_n942), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(G1344gat));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n877), .A2(new_n886), .A3(new_n496), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT57), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n926), .A2(new_n596), .A3(new_n595), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n917), .A2(new_n918), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n670), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n629), .B1(new_n955), .B2(new_n874), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n597), .A2(new_n690), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n931), .B(new_n496), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n933), .A2(new_n688), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n951), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G148gat), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n930), .A2(new_n688), .A3(new_n932), .A4(new_n933), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n336), .A2(KEYINPUT59), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n961), .A2(KEYINPUT59), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n689), .A2(G148gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n939), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n949), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n962), .A2(new_n963), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n960), .B2(G148gat), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n966), .B(KEYINPUT122), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n972), .ZN(G1345gat));
  OAI21_X1  g772(.A(G155gat), .B1(new_n934), .B2(new_n878), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n939), .A2(new_n326), .A3(new_n629), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1346gat));
  OAI21_X1  g775(.A(G162gat), .B1(new_n934), .B2(new_n670), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n908), .A2(new_n327), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n938), .B2(new_n978), .ZN(G1347gat));
  NAND4_X1  g778(.A1(new_n936), .A2(new_n472), .A3(new_n887), .A4(new_n791), .ZN(new_n980));
  INV_X1    g779(.A(G169gat), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n593), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT123), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n695), .A2(new_n472), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT124), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  AOI211_X1 g786(.A(new_n706), .B(new_n987), .C1(new_n894), .C2(new_n895), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n981), .B1(new_n988), .B2(new_n597), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n984), .A2(new_n989), .ZN(G1348gat));
  OR2_X1    g789(.A1(new_n980), .A2(new_n689), .ZN(new_n991));
  INV_X1    g790(.A(G176gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n987), .B1(new_n894), .B2(new_n895), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n706), .A2(new_n249), .A3(new_n689), .ZN(new_n994));
  AOI22_X1  g793(.A1(new_n991), .A2(new_n992), .B1(new_n993), .B2(new_n994), .ZN(G1349gat));
  AOI21_X1  g794(.A(new_n243), .B1(new_n988), .B2(new_n733), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n629), .A2(new_n285), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(KEYINPUT60), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n894), .A2(new_n895), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n1000), .A2(new_n797), .A3(new_n733), .A4(new_n986), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G183gat), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT60), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n1002), .B(new_n1003), .C1(new_n980), .C2(new_n997), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n999), .A2(new_n1004), .ZN(G1350gat));
  NAND3_X1  g804(.A1(new_n993), .A2(new_n797), .A3(new_n669), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n1007));
  AND3_X1   g806(.A1(new_n1006), .A2(new_n1007), .A3(G190gat), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1007), .B1(new_n1006), .B2(G190gat), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n669), .A2(new_n244), .ZN(new_n1010));
  OAI22_X1  g809(.A1(new_n1008), .A2(new_n1009), .B1(new_n980), .B2(new_n1010), .ZN(G1351gat));
  AND2_X1   g810(.A1(new_n951), .A2(new_n958), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n987), .A2(new_n766), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n1014), .A2(new_n361), .A3(new_n714), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n936), .A2(new_n472), .A3(new_n791), .A4(new_n937), .ZN(new_n1016));
  OR2_X1    g815(.A1(new_n1016), .A2(new_n736), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1015), .B1(new_n361), .B2(new_n1017), .ZN(G1352gat));
  OAI21_X1  g817(.A(G204gat), .B1(new_n1014), .B2(new_n689), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n688), .A2(new_n362), .ZN(new_n1020));
  OAI21_X1  g819(.A(KEYINPUT62), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  OR3_X1    g820(.A1(new_n1016), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(G1353gat));
  NAND2_X1  g822(.A1(new_n629), .A2(new_n345), .ZN(new_n1024));
  NOR2_X1   g823(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g824(.A(new_n1025), .B(KEYINPUT125), .Z(new_n1026));
  NAND4_X1  g825(.A1(new_n951), .A2(new_n958), .A3(new_n629), .A4(new_n1013), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1027), .A2(G211gat), .ZN(new_n1028));
  NOR2_X1   g827(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g829(.A(new_n1027), .B(G211gat), .C1(KEYINPUT126), .C2(KEYINPUT63), .ZN(new_n1031));
  NAND2_X1  g830(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1026), .A2(new_n1033), .ZN(G1354gat));
  INV_X1    g833(.A(new_n1014), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n669), .A2(G218gat), .ZN(new_n1036));
  XNOR2_X1  g835(.A(new_n1036), .B(KEYINPUT127), .ZN(new_n1037));
  OR2_X1    g836(.A1(new_n1016), .A2(new_n670), .ZN(new_n1038));
  AOI22_X1  g837(.A1(new_n1035), .A2(new_n1037), .B1(new_n346), .B2(new_n1038), .ZN(G1355gat));
endmodule


