//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n462), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT3), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n461), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n461), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(G100), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n483), .A2(new_n472), .A3(KEYINPUT66), .ZN(new_n484));
  AOI21_X1  g059(.A(KEYINPUT66), .B1(new_n483), .B2(new_n472), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n472), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n471), .A2(G138), .A3(new_n472), .A4(new_n461), .ZN(new_n489));
  INV_X1    g064(.A(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n489), .A2(KEYINPUT4), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT67), .A2(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT67), .A2(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n472), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n472), .A2(G102), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n461), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n493), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT68), .B1(KEYINPUT69), .B2(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT6), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n505), .B1(new_n508), .B2(new_n503), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n502), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n511), .A2(KEYINPUT70), .A3(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT71), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(KEYINPUT72), .A3(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n514), .B1(new_n527), .B2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G89), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n509), .A2(new_n532), .B1(G63), .B2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n509), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n534), .B1(new_n540), .B2(G51), .ZN(G168));
  AOI22_X1  g116(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n507), .ZN(new_n543));
  INV_X1    g118(.A(new_n512), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G90), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n535), .A2(new_n538), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n543), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n518), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n544), .A2(G81), .B1(G651), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n553), .B(KEYINPUT75), .C1(new_n546), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  AOI22_X1  g141(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n507), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n512), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n510), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(new_n572), .A3(G53), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n510), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G51), .ZN(new_n578));
  OAI221_X1 g153(.A(new_n531), .B1(new_n518), .B2(new_n533), .C1(new_n546), .C2(new_n578), .ZN(G286));
  INV_X1    g154(.A(new_n514), .ZN(new_n580));
  INV_X1    g155(.A(new_n528), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT72), .B1(new_n524), .B2(G651), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(G303));
  NAND2_X1  g158(.A1(new_n544), .A2(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n571), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n518), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  INV_X1    g166(.A(G48), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n510), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n512), .A2(KEYINPUT76), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT76), .B1(new_n512), .B2(new_n595), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n544), .A2(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n599), .B1(new_n507), .B2(new_n600), .C1(new_n546), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n536), .A2(KEYINPUT77), .A3(new_n539), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n535), .B2(new_n538), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT10), .B1(new_n544), .B2(G92), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n609), .A2(new_n610), .B1(new_n507), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT78), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n603), .B1(new_n614), .B2(G868), .ZN(G284));
  XOR2_X1   g190(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n576), .B(KEYINPUT80), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n621), .ZN(new_n623));
  MUX2_X1   g198(.A(new_n559), .B(new_n623), .S(G868), .Z(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n479), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n481), .A2(G123), .ZN(new_n628));
  AND2_X1   g203(.A1(G111), .A2(G2105), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G99), .B2(new_n472), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n462), .C2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n490), .A2(new_n474), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT13), .B(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT83), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n652), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(G14), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(new_n654), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n661), .B2(new_n655), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT88), .Z(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT89), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n667), .B(KEYINPUT17), .Z(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n671), .C1(new_n666), .C2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n672), .A3(new_n670), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n665), .A3(new_n667), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(G2096), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n682), .A2(new_n685), .A3(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(G229));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT26), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n479), .A2(G141), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n700), .B(new_n701), .C1(G105), .C2(new_n474), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G129), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT99), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(KEYINPUT100), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT100), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n708), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT101), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G19), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n560), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1341), .Z(new_n719));
  NAND2_X1  g294(.A1(G168), .A2(G16), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT102), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT102), .B1(G16), .B2(G21), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1966), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(G1966), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n711), .B2(new_n713), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n715), .A2(new_n719), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G35), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G162), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2090), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n716), .A2(G20), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT23), .Z(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G299), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1956), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT30), .B(G28), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(G33), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G139), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n743), .B(new_n746), .C1(new_n472), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n742), .B1(new_n748), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n741), .B1(new_n739), .B2(new_n631), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(KEYINPUT24), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(KEYINPUT24), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(KEYINPUT98), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT98), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n476), .B2(new_n739), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n749), .A2(new_n750), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n732), .A2(new_n737), .A3(new_n751), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n614), .B2(G16), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G1348), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G1348), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n739), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  MUX2_X1   g342(.A(G104), .B(G116), .S(G2105), .Z(new_n768));
  AOI22_X1  g343(.A1(new_n481), .A2(G128), .B1(G2104), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n479), .A2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G5), .A2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT103), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G301), .B2(new_n716), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G27), .A2(G29), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G164), .B2(G29), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT104), .B(G2078), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n775), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n761), .A2(new_n764), .A3(new_n765), .A4(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G22), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G166), .B2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(G1971), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n716), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n716), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT33), .B(G1976), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  INV_X1    g373(.A(new_n791), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n792), .A2(KEYINPUT95), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT95), .B1(new_n792), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NOR2_X1   g381(.A1(G25), .A2(G29), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n479), .A2(G131), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT91), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n481), .A2(G119), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n481), .A2(KEYINPUT92), .A3(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G95), .B(G107), .S(G2105), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G2104), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n809), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n807), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  MUX2_X1   g396(.A(G24), .B(G290), .S(G16), .Z(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT93), .B(G1986), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n805), .A2(new_n806), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n805), .A2(new_n828), .A3(new_n806), .A4(new_n825), .ZN(new_n829));
  AOI211_X1 g404(.A(new_n728), .B(new_n786), .C1(new_n827), .C2(new_n829), .ZN(G311));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n829), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n728), .A2(new_n786), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(G150));
  NAND2_X1  g408(.A1(new_n614), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n540), .A2(G55), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n518), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n544), .A2(G93), .B1(G651), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n557), .A3(new_n558), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n555), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n835), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  AOI21_X1  g427(.A(new_n500), .B1(new_n493), .B2(KEYINPUT105), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n490), .A2(new_n492), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n772), .B(new_n859), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n479), .A2(G142), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n481), .A2(G130), .ZN(new_n863));
  MUX2_X1   g438(.A(G106), .B(G118), .S(G2105), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G2104), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n817), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n814), .A2(new_n816), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n809), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT106), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n817), .A2(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n809), .A3(new_n868), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n871), .A2(new_n635), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n635), .B1(new_n871), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n861), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(new_n635), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n871), .A2(new_n635), .A3(new_n875), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n860), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n705), .B(new_n748), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n878), .B2(new_n883), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n487), .B(new_n476), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n631), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n885), .B2(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g469(.A1(new_n841), .A2(G868), .ZN(new_n895));
  XNOR2_X1  g470(.A(G288), .B(KEYINPUT111), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G290), .ZN(new_n897));
  XNOR2_X1  g472(.A(G303), .B(G305), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n613), .B2(G299), .ZN(new_n903));
  OAI211_X1 g478(.A(KEYINPUT107), .B(new_n576), .C1(new_n608), .C2(new_n612), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n613), .A2(G299), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n908), .A3(new_n904), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n907), .A4(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n903), .A2(new_n904), .A3(new_n907), .A4(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT110), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n901), .A2(new_n910), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n623), .B(new_n845), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n623), .B(new_n844), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n911), .A2(new_n907), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n920), .A2(new_n924), .A3(KEYINPUT42), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n910), .A2(new_n901), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n915), .A2(new_n917), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n922), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n900), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n920), .B2(new_n924), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n926), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n899), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n895), .B1(new_n937), .B2(G868), .ZN(G295));
  AOI21_X1  g513(.A(new_n895), .B1(new_n937), .B2(G868), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  NAND3_X1  g515(.A1(G286), .A2(G301), .A3(KEYINPUT112), .ZN(new_n941));
  OAI21_X1  g516(.A(G168), .B1(G301), .B2(KEYINPUT112), .ZN(new_n942));
  AND2_X1   g517(.A1(G301), .A2(KEYINPUT112), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(new_n844), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n922), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n900), .B(new_n946), .C1(new_n918), .C2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n922), .B1(new_n945), .B2(new_n913), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n944), .B(new_n844), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT41), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(new_n910), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n899), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n945), .B1(new_n927), .B2(new_n928), .ZN(new_n956));
  INV_X1    g531(.A(new_n946), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n899), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n953), .A4(new_n947), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n940), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n959), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n953), .A4(new_n947), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n961), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n854), .A2(KEYINPUT105), .A3(new_n855), .ZN(new_n967));
  INV_X1    g542(.A(new_n500), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n493), .A2(KEYINPUT105), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT113), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n853), .B2(new_n858), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n467), .A2(G40), .A3(new_n473), .A4(new_n475), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n705), .B(G1996), .Z(new_n981));
  XNOR2_X1  g556(.A(new_n772), .B(new_n774), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n818), .A2(new_n820), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n818), .A2(new_n820), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(G290), .B(G1986), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n594), .A2(new_n596), .A3(new_n988), .A4(new_n597), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n512), .A2(new_n595), .ZN(new_n990));
  OAI21_X1  g565(.A(G1981), .B1(new_n593), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n973), .B2(new_n978), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n991), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n794), .A2(G1976), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n996), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n996), .B2(new_n1000), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n999), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT50), .B1(new_n859), .B2(new_n966), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT50), .B(new_n966), .C1(new_n493), .C2(new_n500), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n978), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(G2090), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n966), .B1(new_n493), .B2(new_n500), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n977), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1012), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n798), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n995), .B1(new_n1011), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(G166), .B2(new_n995), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1022), .ZN(new_n1024));
  NAND3_X1  g599(.A1(G303), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1006), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT121), .ZN(new_n1028));
  INV_X1    g603(.A(G1966), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1014), .A2(KEYINPUT45), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n1015), .B2(new_n973), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1031), .B2(new_n977), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n758), .B(new_n978), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(G8), .A3(G168), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  NOR3_X1   g613(.A1(G166), .A2(new_n995), .A3(new_n1022), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1024), .B1(G303), .B2(G8), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1023), .A2(new_n1025), .A3(KEYINPUT116), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1013), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(new_n1017), .A3(G1971), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1010), .A2(G2090), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1043), .B(G8), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1006), .B(new_n1048), .C1(new_n1021), .C2(new_n1026), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1028), .A2(new_n1037), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1006), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n859), .B2(new_n966), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1054), .B2(new_n977), .ZN(new_n1055));
  INV_X1    g630(.A(G2090), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT118), .B(new_n978), .C1(new_n973), .C2(new_n1053), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1020), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1020), .A3(KEYINPUT119), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1026), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1035), .B(new_n1051), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1050), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1021), .A2(new_n1006), .A3(new_n1043), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n996), .B(KEYINPUT117), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n999), .A2(G1976), .A3(G288), .ZN(new_n1071));
  INV_X1    g646(.A(new_n989), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT56), .B(G2072), .Z(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n736), .ZN(new_n1080));
  XOR2_X1   g655(.A(new_n576), .B(KEYINPUT57), .Z(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1075), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT118), .B1(new_n1087), .B2(new_n978), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n736), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT123), .A3(new_n1081), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1083), .A2(new_n1085), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1009), .B1(new_n971), .B2(new_n1053), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT122), .B1(new_n1094), .B2(new_n977), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(new_n978), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n973), .A2(new_n774), .A3(new_n978), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(KEYINPUT60), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n614), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n614), .A2(new_n1099), .A3(KEYINPUT60), .A4(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1078), .B(new_n1081), .C1(new_n1079), .C2(new_n736), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1084), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n971), .B2(new_n977), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1076), .B2(G1996), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n560), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT59), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1093), .A2(new_n1108), .A3(new_n1111), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1105), .A2(new_n614), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1083), .A2(new_n1092), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1091), .B2(new_n1081), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n976), .B2(new_n977), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n973), .A2(new_n974), .ZN(new_n1125));
  AOI211_X1 g700(.A(KEYINPUT113), .B(G1384), .C1(new_n853), .C2(new_n858), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1015), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .A3(new_n978), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(G2078), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1013), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1095), .A2(new_n779), .A3(new_n1098), .ZN(new_n1133));
  INV_X1    g708(.A(G2078), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1044), .B2(new_n1017), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1129), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1122), .B1(new_n1137), .B2(G171), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1031), .A2(new_n977), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1130), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1136), .A2(G301), .A3(new_n1133), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT125), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1135), .A2(new_n1129), .B1(new_n1139), .B2(new_n1130), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(G301), .A4(new_n1133), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1133), .ZN(new_n1149));
  OAI21_X1  g724(.A(G171), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1132), .A2(G301), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1122), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1032), .A2(G168), .A3(new_n1033), .ZN(new_n1154));
  AOI21_X1  g729(.A(G168), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT51), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1154), .B(G8), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1154), .A2(G8), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1051), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1147), .A2(new_n1153), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1068), .B(new_n1074), .C1(new_n1121), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1150), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1157), .B(new_n1164), .C1(new_n1158), .C2(new_n1156), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1160), .A2(KEYINPUT126), .A3(new_n1165), .A4(new_n1163), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1168), .A2(new_n1169), .B1(KEYINPUT62), .B2(new_n1159), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n987), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n979), .B1(new_n982), .B2(new_n706), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT127), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n979), .A2(G1996), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT46), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT47), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n981), .A2(new_n982), .ZN(new_n1178));
  OAI22_X1  g753(.A1(new_n1178), .A2(new_n983), .B1(G2067), .B2(new_n772), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n980), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n985), .A2(new_n980), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G290), .A2(G1986), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n980), .A2(KEYINPUT48), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT48), .B1(new_n980), .B2(new_n1182), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1180), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1177), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1171), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g763(.A1(G229), .A2(G227), .A3(new_n457), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n663), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1191), .B1(new_n891), .B2(new_n892), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n1192), .A2(new_n962), .A3(new_n963), .ZN(G308));
  NAND3_X1  g767(.A1(new_n1192), .A2(new_n962), .A3(new_n963), .ZN(G225));
endmodule


