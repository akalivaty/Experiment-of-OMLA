//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT92), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G8gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  AOI21_X1  g004(.A(G1gat), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n204), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT14), .B(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216));
  INV_X1    g015(.A(KEYINPUT91), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n212), .A2(new_n216), .A3(new_n214), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT15), .B1(new_n215), .B2(new_n218), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n222), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n225), .B1(new_n229), .B2(new_n208), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n207), .B(new_n223), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n231), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n225), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n231), .C1(new_n207), .C2(new_n228), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT18), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G169gat), .B(G197gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n245), .B(KEYINPUT12), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n235), .A3(new_n239), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n252));
  AND2_X1   g051(.A1(G211gat), .A2(G218gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(G211gat), .A2(G218gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G197gat), .A2(G204gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n259), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(new_n264), .A3(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n255), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n272));
  AND2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n277), .B(KEYINPUT25), .C1(new_n278), .C2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT66), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n286), .B1(new_n293), .B2(KEYINPUT25), .ZN(new_n294));
  INV_X1    g093(.A(G169gat), .ZN(new_n295));
  INV_X1    g094(.A(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n273), .B1(new_n297), .B2(new_n275), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n281), .B(new_n282), .C1(new_n278), .C2(KEYINPUT66), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n288), .A2(KEYINPUT66), .A3(new_n289), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n272), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n285), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT68), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n308), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT26), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n273), .B1(new_n311), .B2(new_n271), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n288), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT27), .B(G183gat), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT28), .B1(new_n315), .B2(new_n280), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n279), .A2(KEYINPUT27), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G183gat), .ZN(new_n319));
  AND4_X1   g118(.A1(KEYINPUT28), .A2(new_n317), .A3(new_n319), .A4(new_n280), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n305), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n310), .A2(new_n312), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n319), .A3(new_n280), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n280), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n328), .A3(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G226gat), .ZN(new_n331));
  INV_X1    g130(.A(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n304), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n333), .A2(KEYINPUT29), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n288), .A2(new_n289), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n340), .A2(new_n292), .A3(new_n281), .A4(new_n282), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n286), .B(KEYINPUT25), .C1(new_n341), .C2(new_n277), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT67), .B1(new_n301), .B2(new_n302), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n284), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n328), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n337), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n270), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n336), .B1(new_n304), .B2(new_n330), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n345), .A3(new_n333), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n269), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(new_n270), .C1(new_n335), .C2(new_n346), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT30), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n351), .B2(new_n353), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI211_X1 g160(.A(KEYINPUT30), .B(new_n357), .C1(new_n351), .C2(new_n353), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n364));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(G134gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G127gat), .ZN(new_n370));
  INV_X1    g169(.A(G127gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G134gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(KEYINPUT1), .ZN(new_n375));
  INV_X1    g174(.A(G120gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G113gat), .ZN(new_n377));
  INV_X1    g176(.A(G113gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G120gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT76), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n375), .A2(new_n383), .A3(KEYINPUT76), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT74), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G141gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n391), .A3(G148gat), .ZN(new_n392));
  INV_X1    g191(.A(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G141gat), .ZN(new_n394));
  AND2_X1   g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n392), .A2(new_n394), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G155gat), .B(G162gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n388), .A2(G148gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT75), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n395), .A2(new_n397), .ZN(new_n407));
  XNOR2_X1  g206(.A(G141gat), .B(G148gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT2), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n388), .A2(G148gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT74), .B(G141gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(G148gat), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n395), .B1(new_n398), .B2(new_n397), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n406), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(KEYINPUT3), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n394), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n396), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n393), .A2(G141gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n398), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n417), .A2(new_n418), .B1(new_n420), .B2(new_n407), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(KEYINPUT77), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n387), .B(new_n415), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n375), .A2(new_n383), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n375), .A2(new_n383), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n421), .A3(KEYINPUT4), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n428), .A2(new_n429), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n405), .A2(new_n414), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n387), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT79), .B(KEYINPUT5), .C1(new_n439), .C2(new_n433), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n375), .A2(new_n383), .A3(KEYINPUT76), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n405), .B(new_n414), .C1(new_n442), .C2(new_n384), .ZN(new_n443));
  INV_X1    g242(.A(new_n437), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n433), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n434), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n436), .A2(new_n440), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n426), .A2(new_n434), .A3(new_n446), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n364), .B(new_n368), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n451), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n368), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n451), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n451), .A3(new_n368), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n364), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n452), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT87), .B1(new_n363), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n351), .A2(new_n353), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n356), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n358), .ZN(new_n466));
  INV_X1    g265(.A(new_n362), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n368), .B1(new_n453), .B2(new_n454), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n460), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n468), .B(new_n469), .C1(new_n471), .C2(new_n452), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474));
  INV_X1    g273(.A(G50gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT81), .ZN(new_n479));
  INV_X1    g278(.A(G228gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n332), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n421), .A2(new_n416), .A3(new_n422), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n424), .A2(KEYINPUT77), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT29), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(new_n270), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n260), .A2(new_n264), .A3(KEYINPUT82), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n266), .A2(new_n488), .A3(new_n255), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n260), .A2(new_n264), .A3(KEYINPUT82), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(KEYINPUT83), .A3(new_n490), .A4(new_n489), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n422), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n428), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n485), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n490), .A3(new_n489), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT3), .B1(new_n499), .B2(new_n486), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n421), .B1(new_n500), .B2(new_n494), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT84), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n481), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT3), .B1(new_n270), .B2(new_n490), .ZN(new_n504));
  INV_X1    g303(.A(new_n438), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n481), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n485), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n503), .A2(G22gat), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G22gat), .ZN(new_n509));
  OAI22_X1  g308(.A1(new_n501), .A2(KEYINPUT84), .B1(new_n270), .B2(new_n484), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n496), .A2(new_n497), .ZN(new_n511));
  OAI22_X1  g310(.A1(new_n510), .A2(new_n511), .B1(new_n480), .B2(new_n332), .ZN(new_n512));
  INV_X1    g311(.A(new_n507), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n479), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n516), .B(G22gat), .C1(new_n503), .C2(new_n507), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n509), .A3(new_n513), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n478), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n514), .A2(new_n516), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n429), .B1(new_n304), .B2(new_n330), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n328), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT69), .B1(new_n323), .B2(new_n328), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n344), .A2(new_n525), .A3(new_n431), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT64), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT65), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G43gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n531), .B(KEYINPUT32), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n531), .B2(KEYINPUT32), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT33), .B1(new_n527), .B2(new_n530), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT70), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n535), .ZN(new_n541));
  INV_X1    g340(.A(new_n530), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n522), .B2(new_n526), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n545), .A2(new_n546), .A3(new_n538), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n536), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n527), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n529), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT34), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n527), .A2(KEYINPUT34), .A3(new_n530), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555));
  INV_X1    g354(.A(new_n553), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(new_n536), .C1(new_n540), .C2(new_n547), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n521), .A2(new_n554), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n252), .B1(new_n473), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n521), .A2(new_n554), .A3(new_n557), .ZN(new_n560));
  INV_X1    g359(.A(new_n452), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n368), .B1(new_n450), .B2(new_n451), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n460), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n468), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT35), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n560), .C2(new_n564), .ZN(new_n568));
  AND4_X1   g367(.A1(new_n555), .A2(new_n521), .A3(new_n554), .A4(new_n557), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n569), .A2(KEYINPUT88), .A3(new_n472), .A4(new_n463), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n559), .A2(new_n567), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n548), .A2(new_n553), .ZN(new_n572));
  INV_X1    g371(.A(new_n557), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n572), .A2(new_n573), .B1(KEYINPUT71), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n521), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n564), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n356), .B1(new_n464), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n582), .B2(new_n464), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT38), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n348), .A2(new_n349), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n586), .B2(new_n270), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n269), .B1(new_n335), .B2(new_n346), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT38), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n360), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n590), .A3(new_n462), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n430), .A2(new_n432), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n433), .B1(new_n426), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n456), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n439), .A2(new_n433), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT39), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT40), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n363), .A2(new_n458), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n591), .A2(new_n601), .A3(new_n521), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n581), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n251), .B1(new_n571), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n614), .A2(new_n223), .B1(KEYINPUT41), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n228), .B2(new_n614), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G134gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G162gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n618), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(KEYINPUT97), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n619), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G57gat), .B(G64gat), .Z(new_n629));
  XOR2_X1   g428(.A(G71gat), .B(G78gat), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  INV_X1    g431(.A(G71gat), .ZN(new_n633));
  INV_X1    g432(.A(G78gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n629), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n630), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n611), .A2(new_n640), .A3(new_n612), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n611), .B1(new_n640), .B2(new_n612), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT93), .B1(new_n636), .B2(new_n638), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT93), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n651), .B2(new_n613), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n647), .B(new_n613), .C1(new_n653), .C2(new_n648), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n644), .B(new_n646), .C1(new_n652), .C2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n651), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n628), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n644), .B1(new_n652), .B2(new_n655), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n628), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G120gat), .B(G148gat), .Z(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n207), .B1(new_n657), .B2(KEYINPUT21), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT95), .ZN(new_n670));
  NAND2_X1  g469(.A1(G231gat), .A2(G233gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT94), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n670), .B(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT21), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n651), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G127gat), .B(G155gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(G183gat), .B(G211gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n675), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n626), .A2(new_n668), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n604), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n563), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(G1gat), .Z(G1324gat));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n468), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G8gat), .B1(new_n685), .B2(new_n468), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n688), .A2(KEYINPUT101), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n691), .A2(new_n692), .B1(new_n689), .B2(new_n696), .ZN(G1325gat));
  OAI21_X1  g496(.A(G15gat), .B1(new_n685), .B2(new_n579), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n577), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n685), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n521), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n682), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n668), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n626), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n604), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n563), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n213), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n626), .B1(new_n571), .B2(new_n603), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n705), .A2(new_n251), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n715), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n563), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n711), .A2(new_n721), .ZN(G1328gat));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  AOI21_X1  g522(.A(G36gat), .B1(new_n723), .B2(KEYINPUT46), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n707), .A2(new_n363), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n723), .A2(KEYINPUT46), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n720), .B2(new_n468), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  OAI21_X1  g529(.A(G43gat), .B1(new_n720), .B2(new_n579), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n577), .A2(G43gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n604), .A2(new_n706), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT106), .Z(new_n734));
  AOI21_X1  g533(.A(new_n730), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1330gat));
  NAND2_X1  g536(.A1(new_n580), .A2(new_n475), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n707), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n720), .A2(new_n521), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  OAI21_X1  g541(.A(G50gat), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n720), .A2(KEYINPUT109), .A3(new_n521), .ZN(new_n744));
  OAI211_X1 g543(.A(KEYINPUT48), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n741), .B2(new_n475), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n571), .A2(new_n603), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n704), .A2(new_n668), .A3(new_n250), .A4(new_n625), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n708), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g553(.A1(new_n752), .A2(new_n363), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  INV_X1    g558(.A(new_n579), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n633), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n577), .A2(G71gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n752), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n752), .A2(new_n580), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g565(.A1(new_n704), .A2(new_n251), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND4_X1   g568(.A1(KEYINPUT110), .A2(new_n750), .A3(new_n625), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT110), .B1(new_n712), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT111), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n625), .A3(new_n769), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n712), .A2(new_n251), .A3(new_n704), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n768), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n772), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(new_n608), .A3(new_n708), .A4(new_n667), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n668), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n715), .A2(new_n718), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n563), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1336gat));
  NOR3_X1   g585(.A1(new_n668), .A2(G92gat), .A3(new_n468), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT51), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n789), .B2(new_n779), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n777), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n715), .A2(new_n363), .A3(new_n718), .A4(new_n783), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n787), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(new_n794), .B2(G92gat), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n797), .A2(KEYINPUT113), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT113), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(G1337gat));
  NOR3_X1   g600(.A1(new_n577), .A2(G99gat), .A3(new_n668), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n781), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G99gat), .B1(new_n784), .B2(new_n579), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1338gat));
  NOR3_X1   g604(.A1(new_n668), .A2(G106gat), .A3(new_n521), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n791), .B2(new_n792), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n784), .A2(new_n521), .ZN(new_n809));
  INV_X1    g608(.A(G106gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n781), .A2(new_n806), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(new_n659), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n656), .A2(new_n628), .A3(new_n658), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n664), .B1(new_n659), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n820), .A3(KEYINPUT55), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n666), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(new_n818), .B2(new_n820), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(KEYINPUT115), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n825), .B(KEYINPUT55), .C1(new_n818), .C2(new_n820), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n822), .B(new_n829), .C1(new_n824), .C2(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n250), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n230), .A2(new_n231), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n233), .A2(new_n234), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n245), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n249), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n667), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n625), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n625), .A2(new_n835), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n828), .A2(new_n840), .A3(new_n830), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n704), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n683), .A2(new_n250), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT114), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n560), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n363), .A2(new_n563), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n251), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n378), .ZN(G1340gat));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n668), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(new_n376), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n704), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n371), .ZN(G1342gat));
  NAND2_X1  g652(.A1(new_n625), .A2(new_n468), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(G134gat), .A3(new_n563), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT56), .Z(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n847), .B2(new_n626), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1343gat));
  AND2_X1   g658(.A1(new_n579), .A2(new_n846), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n844), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n580), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n822), .A2(new_n250), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n823), .B(KEYINPUT118), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n864), .A2(new_n865), .B1(new_n667), .B2(new_n835), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n625), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n704), .B1(new_n867), .B2(new_n841), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n863), .B(new_n521), .C1(new_n868), .C2(new_n844), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n250), .B(new_n860), .C1(new_n862), .C2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n411), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n861), .A2(new_n708), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n579), .A2(new_n580), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT120), .Z(new_n877));
  AOI21_X1  g676(.A(new_n563), .B1(new_n842), .B2(new_n844), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n251), .A2(G141gat), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n875), .A2(new_n880), .A3(new_n468), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n872), .A2(new_n873), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT58), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n872), .A2(new_n873), .A3(new_n885), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n875), .A2(new_n880), .A3(new_n468), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT59), .B1(new_n888), .B2(new_n668), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n393), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n625), .A2(new_n835), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n866), .A2(new_n625), .B1(new_n891), .B2(new_n827), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n843), .B1(new_n892), .B2(new_n704), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n863), .B1(new_n893), .B2(new_n521), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n896), .B(new_n863), .C1(new_n893), .C2(new_n521), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n863), .B(new_n521), .C1(new_n842), .C2(new_n844), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n860), .A2(new_n667), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT59), .B(G148gat), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n860), .B1(new_n862), .B2(new_n869), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n668), .A2(KEYINPUT59), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n890), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n903), .B2(new_n704), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n704), .A2(G155gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n888), .B2(new_n907), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n903), .B2(new_n626), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n854), .A2(G162gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n875), .A2(new_n880), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1347gat));
  AOI21_X1  g711(.A(new_n708), .B1(new_n842), .B2(new_n844), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n560), .A2(new_n468), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n295), .B1(new_n915), .B2(new_n250), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n914), .B(KEYINPUT123), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n295), .A3(new_n250), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(G1348gat));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n296), .A3(new_n667), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n913), .A2(new_n914), .ZN(new_n923));
  OAI21_X1  g722(.A(G176gat), .B1(new_n923), .B2(new_n668), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1349gat));
  NAND2_X1  g724(.A1(new_n915), .A2(new_n682), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n682), .A2(new_n315), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n926), .A2(G183gat), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n923), .B2(new_n626), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n919), .A2(new_n280), .A3(new_n625), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1351gat));
  NOR2_X1   g733(.A1(new_n876), .A2(new_n468), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT125), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(new_n913), .ZN(new_n937));
  AOI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n250), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n760), .A2(new_n708), .A3(new_n468), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n900), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n250), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  XNOR2_X1  g742(.A(KEYINPUT126), .B(G204gat), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n937), .A2(new_n667), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n667), .B(new_n939), .C1(new_n898), .C2(new_n899), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n947), .B(new_n948), .C1(new_n950), .C2(new_n944), .ZN(G1353gat));
  INV_X1    g750(.A(G211gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n952), .A3(new_n682), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n682), .B(new_n939), .C1(new_n898), .C2(new_n899), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  NAND2_X1  g756(.A1(new_n937), .A2(new_n625), .ZN(new_n958));
  INV_X1    g757(.A(G218gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n626), .A2(new_n959), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n961), .A2(new_n962), .B1(new_n941), .B2(new_n963), .ZN(G1355gat));
endmodule


