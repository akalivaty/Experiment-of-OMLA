//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  OR3_X1    g001(.A1(new_n187), .A2(KEYINPUT66), .A3(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(G137), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(new_n187), .B2(G137), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n188), .B(G131), .C1(new_n190), .C2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(G128), .B(new_n194), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n200), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n187), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n189), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n192), .A2(new_n198), .A3(new_n202), .A4(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n206), .A3(new_n189), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n211), .A2(new_n208), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n199), .A2(new_n200), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT64), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(KEYINPUT30), .B(new_n209), .C1(new_n212), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT2), .A3(G113), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n226), .A2(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n224), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n209), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n216), .A2(new_n218), .A3(new_n222), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n211), .A2(new_n208), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT65), .B1(new_n212), .B2(new_n223), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n234), .B1(new_n241), .B2(KEYINPUT30), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n226), .A2(new_n228), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n229), .A2(new_n230), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n243), .A2(new_n244), .A3(new_n232), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n232), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(new_n209), .C1(new_n212), .C2(new_n223), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n236), .A2(new_n238), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n251), .A2(KEYINPUT68), .A3(new_n209), .A4(new_n247), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n242), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n255), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT29), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n239), .A2(new_n240), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n247), .B1(new_n263), .B2(new_n209), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n250), .A2(new_n252), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT28), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n248), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n260), .B(KEYINPUT71), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(KEYINPUT72), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n268), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n250), .B(new_n252), .C1(new_n241), .C2(new_n247), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(KEYINPUT28), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT72), .B1(new_n275), .B2(new_n270), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n209), .B1(new_n212), .B2(new_n223), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n233), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n250), .A2(new_n252), .A3(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n279), .B(new_n273), .C1(new_n282), .C2(KEYINPUT28), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n278), .B1(new_n283), .B2(G902), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n268), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT73), .B(new_n285), .C1(new_n287), .C2(new_n279), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n277), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n224), .A2(new_n233), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n212), .A2(new_n223), .A3(KEYINPUT65), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n209), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n250), .A2(new_n252), .A3(new_n260), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT70), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n242), .A2(new_n253), .A3(new_n300), .A4(new_n260), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n242), .A2(new_n253), .A3(new_n303), .A4(new_n260), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n275), .B2(new_n270), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n291), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n301), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n295), .A2(new_n233), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n267), .B1(new_n310), .B2(new_n253), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n269), .B1(new_n311), .B2(new_n273), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n312), .A3(new_n304), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n290), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G140), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n317), .A3(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G146), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n316), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n196), .B1(new_n326), .B2(new_n317), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(KEYINPUT75), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(G146), .B1(new_n328), .B2(new_n323), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .B1(new_n317), .B2(new_n326), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT76), .B1(new_n335), .B2(G146), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(G128), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT74), .A3(G110), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT74), .B1(new_n343), .B2(G110), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n201), .A2(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n342), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT24), .B(G110), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(new_n344), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n327), .A2(new_n328), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n334), .B2(new_n196), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n354), .A2(new_n318), .A3(new_n320), .A4(new_n196), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n358));
  INV_X1    g172(.A(G110), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n358), .A2(new_n359), .B1(new_n347), .B2(new_n348), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n352), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n356), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n334), .A2(new_n196), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n347), .A2(new_n348), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n343), .B2(G110), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT78), .A4(new_n353), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n351), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G953), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G221), .A3(G234), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT79), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G137), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n351), .A2(new_n369), .A3(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G234), .ZN(new_n380));
  OAI21_X1  g194(.A(G217), .B1(new_n380), .B2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n285), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n382), .B(KEYINPUT81), .Z(new_n383));
  NOR2_X1   g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n285), .A3(new_n378), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT80), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n381), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n315), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G214), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(G107), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G104), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(G104), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(KEYINPUT3), .C1(new_n396), .C2(G107), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n398), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(G101), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n398), .B(new_n407), .C1(new_n401), .C2(new_n403), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT82), .B1(new_n397), .B2(new_n395), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n402), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n407), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n233), .B(new_n406), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n396), .A2(G107), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n410), .B2(new_n402), .ZN(new_n416));
  XNOR2_X1  g230(.A(G104), .B(G107), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT84), .B1(new_n417), .B2(new_n407), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(G101), .C1(new_n397), .C2(new_n394), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n416), .A2(new_n407), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n245), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n339), .A2(G116), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n423), .B(G113), .C1(KEYINPUT5), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n413), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n413), .A2(new_n426), .A3(new_n428), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n198), .A2(new_n202), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n319), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n236), .B2(new_n319), .ZN(new_n435));
  INV_X1    g249(.A(G224), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G953), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n428), .B1(new_n413), .B2(new_n426), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n432), .B(new_n438), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(new_n436), .B2(G953), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n428), .B(KEYINPUT8), .Z(new_n447));
  NAND2_X1  g261(.A1(new_n422), .A2(new_n425), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n418), .A2(new_n420), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n408), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n447), .B1(new_n426), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n435), .A2(new_n445), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n446), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(G902), .B1(new_n454), .B2(new_n431), .ZN(new_n455));
  OAI21_X1  g269(.A(G210), .B1(G237), .B2(G902), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n444), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n444), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n392), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n396), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n365), .B1(new_n196), .B2(new_n334), .ZN(new_n463));
  INV_X1    g277(.A(G237), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n371), .A3(G214), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(G143), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n193), .A2(KEYINPUT87), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G214), .A3(new_n256), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT18), .A2(G131), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n469), .B1(G214), .B2(new_n256), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n465), .A2(new_n467), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n470), .A3(new_n207), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n334), .B(KEYINPUT19), .Z(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(new_n353), .C1(new_n480), .C2(G146), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n462), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n463), .A2(new_n473), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n484), .A3(new_n478), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n471), .A2(KEYINPUT17), .A3(G131), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(KEYINPUT88), .B2(new_n337), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n330), .A2(new_n336), .A3(new_n489), .A4(new_n333), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n483), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n482), .B1(new_n491), .B2(new_n462), .ZN(new_n492));
  NOR2_X1   g306(.A1(G475), .A2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT20), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n327), .A2(KEYINPUT75), .A3(new_n328), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT75), .B1(new_n327), .B2(new_n328), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n496), .A2(new_n497), .B1(new_n332), .B2(new_n331), .ZN(new_n498));
  INV_X1    g312(.A(new_n333), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT88), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n487), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n490), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n462), .A3(new_n474), .ZN(new_n503));
  INV_X1    g317(.A(new_n482), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n493), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n474), .ZN(new_n509));
  INV_X1    g323(.A(new_n462), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n511), .B2(new_n503), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT90), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n502), .A2(new_n462), .A3(new_n474), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n462), .B1(new_n502), .B2(new_n474), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT90), .B(new_n285), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT89), .B(G475), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n508), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G116), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT14), .A3(G122), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(G122), .ZN(new_n523));
  INV_X1    g337(.A(G122), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G116), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(G107), .B(new_n522), .C1(new_n526), .C2(KEYINPUT14), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n525), .A3(new_n393), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n201), .A2(G143), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n201), .A2(G143), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n187), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n187), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n527), .B(new_n528), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n528), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n393), .B1(new_n523), .B2(new_n525), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT91), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n526), .A2(G107), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n528), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n541), .A3(new_n532), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n201), .B2(G143), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n193), .A2(KEYINPUT13), .A3(G128), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n531), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n546), .A2(new_n547), .A3(G134), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n546), .B2(G134), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n535), .B1(new_n542), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT9), .B(G234), .ZN(new_n552));
  INV_X1    g366(.A(G217), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(G953), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n535), .B(new_n554), .C1(new_n542), .C2(new_n550), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n285), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT93), .B1(new_n558), .B2(new_n285), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n564), .B(G902), .C1(new_n556), .C2(new_n557), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n562), .B1(new_n566), .B2(new_n561), .ZN(new_n567));
  NAND2_X1  g381(.A1(G234), .A2(G237), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(G952), .A3(new_n371), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT94), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT21), .B(G898), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n568), .A2(G902), .A3(G953), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n520), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n392), .C1(new_n457), .C2(new_n458), .ZN(new_n579));
  INV_X1    g393(.A(G469), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n450), .A2(new_n433), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n198), .A2(new_n202), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n408), .B2(new_n449), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n238), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT12), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n236), .B(new_n406), .C1(new_n409), .C2(new_n412), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n421), .B2(new_n582), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n582), .A2(new_n408), .A3(new_n449), .A4(new_n587), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n212), .B(new_n586), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(G110), .B(G140), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n371), .A2(G227), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n238), .C1(new_n581), .C2(new_n583), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n585), .A2(new_n591), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n238), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n595), .B1(new_n601), .B2(new_n591), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n580), .B(new_n285), .C1(new_n599), .C2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n580), .A2(new_n285), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n585), .A2(new_n591), .A3(new_n597), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n594), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n601), .A2(new_n591), .A3(new_n595), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(G469), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G221), .B1(new_n552), .B2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n460), .A2(new_n577), .A3(new_n579), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n391), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n407), .ZN(G3));
  AND3_X1   g430(.A1(new_n390), .A2(new_n610), .A3(new_n611), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n313), .A2(new_n285), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(G472), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n266), .A2(new_n268), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n297), .A2(new_n298), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n621), .A2(new_n269), .B1(new_n622), .B2(new_n303), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n623), .B2(new_n309), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT95), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n617), .A2(new_n306), .A3(new_n620), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n566), .A2(new_n560), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n558), .B(KEYINPUT33), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n560), .A2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n520), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n392), .B(new_n575), .C1(new_n457), .C2(new_n458), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  OAI21_X1  g453(.A(new_n285), .B1(new_n514), .B2(new_n515), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT90), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n518), .A3(new_n516), .ZN(new_n643));
  INV_X1    g457(.A(new_n563), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n558), .A2(KEYINPUT93), .A3(new_n285), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n561), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n562), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n495), .A2(new_n649), .A3(new_n507), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT20), .B(new_n494), .C1(new_n503), .C2(new_n504), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT96), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n643), .A2(new_n648), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n635), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n628), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n376), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n370), .B(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n383), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n388), .B2(new_n389), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n620), .A2(new_n626), .A3(new_n306), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n614), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT37), .B(G110), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  NOR2_X1   g483(.A1(new_n459), .A2(new_n612), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n315), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n573), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n570), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n672), .B1(new_n653), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n519), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n567), .B1(new_n677), .B2(new_n642), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n507), .A2(new_n649), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n506), .B1(new_n505), .B2(new_n493), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n651), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n679), .B1(new_n681), .B2(new_n649), .ZN(new_n682));
  INV_X1    g496(.A(new_n675), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n678), .A2(new_n682), .A3(KEYINPUT99), .A4(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(new_n458), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n444), .A2(new_n455), .A3(new_n456), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n392), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n665), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n675), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n613), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n520), .A2(new_n648), .ZN(new_n699));
  INV_X1    g513(.A(new_n291), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n307), .B(new_n700), .C1(new_n623), .C2(new_n309), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT32), .B1(new_n313), .B2(new_n291), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n269), .A2(new_n282), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n299), .A2(new_n301), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(KEYINPUT101), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(KEYINPUT101), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n699), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n694), .A2(new_n697), .A3(new_n698), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n643), .A2(new_n508), .B1(new_n629), .B2(new_n632), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n683), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n712), .A2(new_n520), .A3(new_n633), .A4(new_n683), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n664), .B1(new_n703), .B2(new_n290), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n670), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  INV_X1    g533(.A(new_n591), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT10), .B1(new_n450), .B2(new_n433), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n589), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n212), .B1(new_n722), .B2(new_n586), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n594), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n598), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n580), .B1(new_n725), .B2(new_n285), .ZN(new_n726));
  AOI211_X1 g540(.A(G469), .B(G902), .C1(new_n724), .C2(new_n598), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT103), .B1(new_n728), .B2(new_n611), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  INV_X1    g544(.A(new_n611), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n726), .A2(new_n727), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n315), .A3(new_n390), .A4(new_n636), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n735));
  INV_X1    g549(.A(new_n390), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n703), .B2(new_n290), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n636), .A4(new_n733), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND4_X1  g556(.A1(new_n733), .A2(new_n654), .A3(new_n315), .A4(new_n390), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NAND3_X1  g558(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n611), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n285), .B1(new_n599), .B2(new_n602), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n611), .A3(new_n603), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n730), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n693), .B1(new_n688), .B2(new_n689), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n315), .A3(new_n577), .A4(new_n665), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  AOI21_X1  g567(.A(new_n625), .B1(new_n313), .B2(new_n285), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n287), .A2(new_n269), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n304), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n700), .B1(new_n757), .B2(new_n309), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n736), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n699), .A2(new_n459), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n733), .A3(new_n575), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NAND3_X1  g576(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n618), .A2(G472), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n291), .B1(new_n302), .B2(new_n756), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n665), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n716), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  XNOR2_X1  g583(.A(new_n702), .B(KEYINPUT107), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n290), .A2(new_n314), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n390), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n520), .A2(new_n633), .A3(new_n683), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT102), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n606), .A2(new_n775), .A3(new_n594), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n608), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n775), .B1(new_n606), .B2(new_n594), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n580), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n603), .A2(new_n605), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n611), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n688), .A2(new_n392), .A3(new_n689), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n713), .A2(new_n712), .A3(new_n683), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n774), .A2(new_n783), .A3(new_n784), .A4(KEYINPUT42), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n772), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n315), .A2(new_n783), .A3(new_n390), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n774), .A2(new_n784), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT106), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n792), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n786), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n207), .ZN(G33));
  NAND4_X1  g609(.A1(new_n685), .A2(KEYINPUT108), .A3(new_n737), .A4(new_n783), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n676), .A2(new_n684), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n788), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G134), .ZN(G36));
  NAND2_X1  g615(.A1(new_n607), .A2(KEYINPUT105), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT45), .A3(new_n608), .A4(new_n776), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n607), .A2(new_n608), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n803), .B(G469), .C1(KEYINPUT45), .C2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n605), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(KEYINPUT46), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n603), .B1(new_n806), .B2(KEYINPUT46), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n611), .B(new_n695), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n643), .A2(new_n633), .A3(new_n508), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT43), .Z(new_n812));
  NAND3_X1  g626(.A1(new_n620), .A2(new_n626), .A3(new_n306), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n665), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n809), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n810), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n782), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT109), .B(G137), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G39));
  OAI21_X1  g634(.A(new_n611), .B1(new_n807), .B2(new_n808), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT47), .Z(new_n822));
  NOR4_X1   g636(.A1(new_n789), .A2(new_n315), .A3(new_n390), .A4(new_n782), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  NAND3_X1  g639(.A1(new_n390), .A2(new_n392), .A3(new_n611), .ZN(new_n826));
  INV_X1    g640(.A(new_n728), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n811), .B(new_n826), .C1(KEYINPUT49), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT110), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n703), .A2(new_n708), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT111), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n829), .A2(new_n692), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n812), .A2(new_n571), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n759), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n692), .A2(new_n733), .A3(new_n693), .ZN(new_n837));
  OR4_X1    g651(.A1(KEYINPUT116), .A2(new_n836), .A3(KEYINPUT50), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n729), .A2(new_n732), .A3(new_n782), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(new_n766), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n831), .A2(new_n390), .A3(new_n571), .A4(new_n841), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n844), .A2(new_n520), .A3(new_n633), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n840), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n821), .B(KEYINPUT47), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n728), .A2(new_n731), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n782), .B(new_n836), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT117), .B1(new_n850), .B2(KEYINPUT51), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n844), .A2(new_n634), .ZN(new_n852));
  INV_X1    g666(.A(G952), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(new_n853), .A3(G953), .ZN(new_n854));
  INV_X1    g668(.A(new_n772), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n835), .A3(new_n841), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  OAI221_X1 g672(.A(new_n854), .B1(new_n763), .B2(new_n836), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n850), .B2(KEYINPUT51), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n861), .B(new_n862), .C1(new_n846), .C2(new_n849), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n851), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n614), .B1(new_n391), .B2(new_n666), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n643), .A2(new_n508), .A3(new_n648), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n634), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n460), .A3(new_n579), .A4(new_n575), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n627), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n643), .A2(new_n567), .A3(new_n683), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n650), .A2(new_n652), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n664), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n315), .A2(new_n874), .A3(new_n613), .ZN(new_n875));
  AOI21_X1  g689(.A(G902), .B1(new_n724), .B2(new_n598), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n604), .B1(new_n876), .B2(new_n580), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n802), .A2(G469), .A3(new_n608), .A4(new_n776), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n731), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n764), .A2(new_n665), .A3(new_n765), .A4(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n875), .B1(new_n789), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n782), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n800), .A2(new_n871), .A3(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n772), .A2(new_n785), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n716), .A2(new_n737), .A3(new_n783), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n792), .B1(new_n886), .B2(new_n787), .ZN(new_n887));
  INV_X1    g701(.A(new_n793), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n671), .A2(new_n685), .B1(new_n767), .B2(new_n716), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n664), .A2(new_n683), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT113), .B1(new_n892), .B2(new_n781), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n879), .A2(new_n894), .A3(new_n664), .A4(new_n683), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n709), .A3(new_n750), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n890), .A2(new_n891), .A3(new_n718), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n686), .A2(new_n718), .A3(new_n897), .A4(new_n768), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT52), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n884), .A2(new_n889), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n735), .A2(new_n739), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n752), .A2(new_n743), .A3(new_n761), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT112), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n752), .A2(new_n743), .A3(new_n761), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT112), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n740), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n865), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n740), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n905), .B2(new_n740), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n900), .A2(new_n898), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n800), .A2(new_n871), .A3(new_n883), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n794), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n865), .B1(new_n890), .B2(new_n891), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n912), .A2(new_n913), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT54), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT114), .B1(new_n902), .B2(new_n903), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT114), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n905), .A2(new_n921), .A3(new_n740), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n890), .A2(new_n891), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n865), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n913), .A2(new_n923), .A3(new_n915), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n909), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n919), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n864), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(G952), .A2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n834), .B1(new_n930), .B2(new_n931), .ZN(G75));
  NAND2_X1  g746(.A1(new_n853), .A2(G953), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT119), .Z(new_n934));
  AOI21_X1  g748(.A(new_n285), .B1(new_n909), .B2(new_n926), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(G210), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n438), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n939), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT118), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT118), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n936), .A2(new_n943), .A3(new_n939), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(G51));
  INV_X1    g759(.A(new_n934), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n725), .B(KEYINPUT120), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n909), .A2(new_n927), .A3(new_n926), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n927), .B1(new_n909), .B2(new_n926), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n604), .B(KEYINPUT57), .Z(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n935), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(new_n805), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n946), .B1(new_n952), .B2(new_n954), .ZN(G54));
  NAND3_X1  g769(.A1(new_n935), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n956), .A2(KEYINPUT121), .A3(new_n492), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n934), .B1(new_n956), .B2(new_n492), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT121), .B1(new_n956), .B2(new_n492), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n630), .B1(new_n929), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n630), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n963), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n948), .B2(new_n949), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n934), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n961), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT54), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n909), .B2(new_n917), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n948), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n966), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(KEYINPUT122), .A3(new_n934), .A4(new_n968), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n909), .B2(new_n926), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n379), .B(KEYINPUT123), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n661), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n934), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n934), .A4(new_n982), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G66));
  INV_X1    g801(.A(new_n572), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n371), .B1(new_n988), .B2(G224), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n912), .A2(new_n871), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n371), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n937), .B1(G898), .B2(new_n371), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n991), .B(new_n992), .Z(G69));
  AND2_X1   g807(.A1(new_n890), .A2(new_n718), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n855), .A2(new_n760), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n994), .B(new_n800), .C1(new_n809), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(new_n794), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n822), .A2(new_n823), .B1(new_n817), .B2(new_n815), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n371), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n224), .B1(new_n241), .B2(KEYINPUT30), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(new_n480), .Z(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(G900), .B2(G953), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n371), .B1(G227), .B2(G900), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n1000), .A2(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n696), .A2(new_n782), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n737), .A2(new_n868), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n994), .A2(new_n710), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1010), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1014));
  AOI21_X1  g828(.A(KEYINPUT124), .B1(new_n1010), .B2(KEYINPUT62), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1013), .B(new_n998), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n371), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n1002), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1005), .A2(new_n1004), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(G72));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(new_n1016), .B2(new_n990), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n260), .A3(new_n254), .ZN(new_n1025));
  INV_X1    g839(.A(new_n254), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1026), .A2(new_n260), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1028), .A2(KEYINPUT127), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n299), .B(new_n301), .C1(new_n1028), .C2(KEYINPUT127), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n918), .B(new_n1023), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1023), .ZN(new_n1033));
  INV_X1    g847(.A(new_n990), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1033), .B1(new_n999), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1026), .A2(new_n261), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n934), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT126), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1039), .B(new_n934), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1032), .B1(new_n1038), .B2(new_n1040), .ZN(G57));
endmodule


