//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  OR3_X1    g0018(.A1(new_n217), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n215), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT64), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(G1698), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n254), .B1(new_n255), .B2(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n248), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(new_n265), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n262), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(G226), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n210), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(G20), .B2(new_n203), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n218), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n209), .A2(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G50), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G50), .B2(new_n284), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n272), .A2(G169), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(KEYINPUT65), .B1(new_n291), .B2(new_n272), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(KEYINPUT65), .B2(new_n290), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n283), .A2(new_n289), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT9), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G190), .B2(new_n272), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT66), .B(G200), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n271), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT67), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n296), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n296), .B2(new_n301), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n293), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n277), .A2(new_n202), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n274), .A2(new_n255), .B1(new_n210), .B2(G68), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n281), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT11), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT69), .B1(new_n284), .B2(G68), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT12), .Z(new_n312));
  NAND3_X1  g0112(.A1(new_n286), .A2(G68), .A3(new_n287), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n308), .A2(new_n309), .ZN(new_n314));
  AND4_X1   g0114(.A1(new_n310), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n266), .B1(new_n268), .B2(new_n222), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  INV_X1    g0119(.A(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n256), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G226), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n318), .B(new_n319), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n317), .B1(new_n323), .B2(new_n260), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n326), .B(G179), .C1(new_n327), .C2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n324), .A2(new_n327), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(G179), .A4(new_n326), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n323), .A2(new_n260), .ZN(new_n334));
  INV_X1    g0134(.A(new_n317), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n334), .A2(new_n325), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n324), .A2(new_n325), .ZN(new_n337));
  OAI21_X1  g0137(.A(G169), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT14), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(G169), .C1(new_n336), .C2(new_n337), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n316), .B1(new_n333), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n330), .A2(G190), .A3(new_n326), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n315), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n336), .A2(new_n337), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(G200), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n273), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n351), .B1(new_n274), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n281), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n286), .A2(G77), .A3(new_n287), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(G77), .C2(new_n284), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n258), .A2(new_n222), .B1(new_n206), .B2(new_n256), .ZN(new_n360));
  INV_X1    g0160(.A(G232), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n252), .A2(new_n361), .A3(G1698), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n260), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n267), .B1(G244), .B2(new_n269), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n359), .B1(G169), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n365), .A2(G179), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n359), .B1(G190), .B2(new_n366), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n298), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n305), .A2(new_n349), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n252), .B2(new_n210), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n377), .B(G20), .C1(new_n249), .C2(new_n251), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n221), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n276), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n377), .B1(new_n256), .B2(G20), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n250), .A2(G33), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT7), .B(new_n210), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n221), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n387), .B1(new_n392), .B2(new_n384), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n393), .A3(new_n281), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n386), .A2(new_n393), .A3(KEYINPUT71), .A4(new_n281), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n286), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n350), .A2(new_n287), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(new_n284), .B2(new_n350), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n256), .A2(G226), .A3(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT72), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n256), .A2(new_n407), .A3(G226), .A4(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n253), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n265), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n266), .B1(new_n268), .B2(new_n361), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n412), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n321), .A2(new_n257), .B1(new_n248), .B2(new_n223), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n408), .B2(new_n406), .ZN(new_n416));
  OAI211_X1 g0216(.A(G179), .B(new_n414), .C1(new_n416), .C2(new_n265), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n403), .A2(new_n404), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n401), .B1(new_n396), .B2(new_n397), .ZN(new_n420));
  INV_X1    g0220(.A(new_n418), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT18), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT73), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n411), .B2(new_n412), .ZN(new_n426));
  INV_X1    g0226(.A(G190), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n414), .C1(new_n416), .C2(new_n265), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AND4_X1   g0229(.A1(KEYINPUT17), .A2(new_n398), .A3(new_n402), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT17), .B1(new_n420), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n424), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n379), .A2(new_n385), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n282), .B1(new_n433), .B2(new_n387), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT71), .B1(new_n434), .B2(new_n386), .ZN(new_n435));
  INV_X1    g0235(.A(new_n397), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n402), .B(new_n429), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n420), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n423), .B1(new_n432), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n375), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  INV_X1    g0244(.A(G169), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n260), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n447), .ZN(new_n450));
  INV_X1    g0250(.A(G274), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n260), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n449), .A2(G270), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n249), .A2(new_n251), .A3(G264), .A4(G1698), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n249), .A2(new_n251), .A3(G257), .A4(new_n320), .ZN(new_n455));
  INV_X1    g0255(.A(G303), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n256), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n260), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n445), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n448), .A2(new_n447), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G270), .A3(new_n265), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n448), .A2(new_n265), .A3(G274), .A4(new_n447), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n260), .B2(new_n457), .ZN(new_n464));
  AOI22_X1  g0264(.A1(KEYINPUT21), .A2(new_n459), .B1(new_n464), .B2(G179), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n280), .A2(new_n218), .B1(G20), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT20), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n285), .A2(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n209), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n284), .A2(new_n474), .A3(new_n218), .A4(new_n280), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(G116), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT78), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n467), .A2(new_n469), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n284), .A2(new_n466), .ZN(new_n484));
  INV_X1    g0284(.A(new_n475), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n466), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT78), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n444), .B1(new_n465), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n457), .A2(new_n260), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT21), .B(G169), .C1(new_n490), .C2(new_n463), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n453), .A2(G179), .A3(new_n458), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n477), .B1(new_n472), .B2(new_n476), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n483), .A2(KEYINPUT78), .A3(new_n486), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n496), .ZN(new_n497));
  AOI211_X1 g0297(.A(KEYINPUT80), .B(KEYINPUT21), .C1(new_n496), .C2(new_n459), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n459), .B1(new_n478), .B2(new_n487), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n489), .B(new_n497), .C1(new_n498), .C2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n488), .B(KEYINPUT81), .C1(new_n425), .C2(new_n464), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n464), .A2(new_n425), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(new_n496), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n464), .A2(G190), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n504), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n460), .A2(G257), .A3(new_n265), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n462), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n249), .A2(new_n251), .A3(G244), .A4(new_n320), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n468), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n260), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n512), .A2(new_n521), .A3(new_n462), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n514), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n525), .A2(new_n205), .A3(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G97), .B(G107), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n528), .A2(new_n210), .B1(new_n255), .B2(new_n277), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n206), .B1(new_n388), .B2(new_n391), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n281), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n485), .A2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n285), .A2(new_n205), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n513), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n520), .A3(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n524), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n520), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n445), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n531), .A2(new_n534), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n514), .A2(new_n291), .A3(new_n520), .A4(new_n522), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(G20), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT84), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT85), .B1(new_n206), .B2(G20), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(KEYINPUT23), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n210), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n550), .A2(new_n552), .B1(new_n553), .B2(KEYINPUT84), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n256), .A2(new_n557), .A3(new_n210), .A4(G87), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n249), .A2(new_n251), .A3(new_n210), .A4(G87), .ZN(new_n559));
  XOR2_X1   g0359(.A(KEYINPUT82), .B(KEYINPUT22), .Z(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n555), .A2(new_n556), .A3(new_n558), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(new_n561), .A3(new_n549), .A4(new_n554), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT83), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n562), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n281), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT25), .B1(new_n285), .B2(new_n206), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n285), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n570), .A2(new_n571), .B1(G107), .B2(new_n485), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G294), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(new_n320), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n260), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n449), .A2(G264), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n462), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n425), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n580), .A2(KEYINPUT86), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(KEYINPUT86), .C1(G190), .C2(new_n579), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n568), .A2(new_n572), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n260), .A2(new_n224), .A3(new_n447), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n265), .A2(G274), .ZN(new_n586));
  INV_X1    g0386(.A(new_n447), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n265), .A2(KEYINPUT75), .A3(G274), .A4(new_n447), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n256), .A2(G238), .A3(new_n320), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n256), .A2(G244), .A3(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n545), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n260), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(G190), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n590), .A2(new_n594), .A3(KEYINPUT77), .A4(G190), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n256), .A2(new_n210), .A3(G68), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n210), .B1(new_n319), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G87), .B2(new_n207), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT76), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n604), .A2(new_n605), .A3(new_n601), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n604), .B2(new_n601), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n600), .B(new_n603), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n281), .B1(new_n285), .B2(new_n355), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n485), .A2(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n297), .B1(new_n590), .B2(new_n594), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n590), .A2(new_n594), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n485), .A2(new_n354), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n445), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n590), .A2(new_n291), .A3(new_n594), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n599), .A2(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n544), .A2(new_n583), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n579), .A2(new_n445), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G179), .B2(new_n579), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n562), .A2(new_n564), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT24), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n282), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n572), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n443), .A2(new_n511), .A3(new_n629), .ZN(G372));
  OAI21_X1  g0430(.A(new_n343), .B1(new_n347), .B2(new_n370), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT73), .B1(new_n439), .B2(new_n440), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n439), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n423), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n304), .B2(new_n303), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n293), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n621), .B1(new_n568), .B2(new_n572), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n500), .A2(new_n501), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT80), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n500), .A2(new_n499), .A3(new_n501), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n488), .B2(new_n465), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n619), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n616), .A2(new_n617), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT87), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n543), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n618), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n618), .A2(KEYINPUT26), .A3(new_n650), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT88), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n647), .B(KEYINPUT87), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n618), .A2(KEYINPUT26), .A3(new_n650), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT26), .B1(new_n618), .B2(new_n650), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n656), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n646), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n639), .B1(new_n443), .B2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n488), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n645), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n511), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n671), .B1(new_n626), .B2(new_n627), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n640), .B1(new_n678), .B2(new_n583), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n628), .A2(new_n671), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT89), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n583), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n628), .ZN(new_n683));
  INV_X1    g0483(.A(new_n680), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT89), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n677), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n496), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT79), .B1(new_n493), .B2(new_n496), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n671), .B1(new_n690), .B2(new_n644), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n686), .A2(new_n681), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n684), .A3(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n213), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n217), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n661), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n671), .B1(new_n703), .B2(new_n646), .ZN(new_n704));
  XNOR2_X1  g0504(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n544), .A2(new_n583), .A3(new_n618), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n690), .A2(new_n628), .A3(new_n644), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT91), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n690), .A2(new_n628), .A3(new_n644), .A4(KEYINPUT91), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n701), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n709), .B1(new_n715), .B2(new_n671), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n712), .B1(new_n503), .B2(new_n640), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n619), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n655), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT92), .A3(new_n672), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n708), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  AOI211_X1 g0523(.A(KEYINPUT93), .B(new_n723), .C1(new_n716), .C2(new_n720), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n707), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n510), .A2(new_n619), .A3(new_n628), .A4(new_n672), .ZN(new_n726));
  INV_X1    g0526(.A(new_n539), .ZN(new_n727));
  INV_X1    g0527(.A(new_n614), .ZN(new_n728));
  INV_X1    g0528(.A(new_n492), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n576), .A2(new_n260), .B1(G264), .B2(new_n449), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n728), .A2(G179), .A3(new_n464), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n579), .A3(new_n523), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(new_n732), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n671), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n726), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n725), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n700), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(G13), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n209), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n695), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n675), .A2(G330), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n677), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n210), .A2(new_n291), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OR3_X1    g0555(.A1(new_n755), .A2(KEYINPUT97), .A3(new_n425), .ZN(new_n756));
  OAI21_X1  g0556(.A(KEYINPUT97), .B1(new_n755), .B2(new_n425), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n427), .A3(new_n757), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT100), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT100), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n756), .A2(G190), .A3(new_n757), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G326), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n755), .A2(new_n427), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n210), .A2(G179), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n767), .A2(G322), .B1(G329), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n754), .A2(new_n769), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n772), .B(new_n252), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n427), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n210), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n775), .B1(G294), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n298), .A2(new_n768), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n427), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G283), .A2(new_n781), .B1(new_n782), .B2(G303), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n763), .A2(new_n766), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n774), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n781), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n255), .B1(new_n790), .B2(new_n206), .ZN(new_n791));
  INV_X1    g0591(.A(new_n782), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n223), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n778), .A2(G97), .ZN(new_n795));
  INV_X1    g0595(.A(new_n767), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n256), .B(new_n795), .C1(new_n796), .C2(new_n380), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT98), .B(G159), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n770), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n800));
  XNOR2_X1  g0600(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n794), .B(new_n802), .C1(new_n202), .C2(new_n764), .ZN(new_n803));
  INV_X1    g0603(.A(new_n761), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n221), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n784), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n218), .B1(G20), .B2(new_n445), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n746), .A2(new_n248), .A3(KEYINPUT95), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT95), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(G13), .B2(G33), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n807), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n213), .A2(new_n252), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT94), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n246), .A2(G45), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G45), .C2(new_n217), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n694), .A2(new_n252), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G355), .B1(new_n466), .B2(new_n694), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n806), .A2(new_n807), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n813), .B(KEYINPUT101), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n675), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n750), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n753), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT102), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n359), .A2(new_n671), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n373), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n370), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n369), .A2(new_n672), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n704), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n750), .B1(new_n835), .B2(new_n743), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n743), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n781), .A2(G68), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n252), .B1(new_n771), .B2(G132), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n838), .B(new_n839), .C1(new_n380), .C2(new_n777), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n767), .A2(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n764), .B2(new_n842), .C1(new_n789), .C2(new_n798), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G150), .B2(new_n761), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n840), .B(new_n845), .C1(G50), .C2(new_n782), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n781), .A2(G87), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n792), .B2(new_n206), .C1(new_n789), .C2(new_n466), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n765), .A2(G303), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n767), .A2(G294), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n256), .B1(new_n771), .B2(G311), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n849), .A2(new_n795), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n848), .B(new_n852), .C1(G283), .C2(new_n761), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n807), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n811), .A2(new_n807), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n750), .B1(G77), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT103), .Z(new_n858));
  OAI211_X1 g0658(.A(new_n854), .B(new_n858), .C1(new_n812), .C2(new_n834), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n837), .A2(new_n859), .ZN(G384));
  NOR3_X1   g0660(.A1(new_n218), .A2(new_n210), .A3(new_n466), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n528), .B(KEYINPUT104), .Z(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OR3_X1    g0667(.A1(new_n217), .A2(new_n255), .A3(new_n381), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n202), .A2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n209), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n343), .A2(new_n671), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n635), .B1(new_n633), .B2(new_n632), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n401), .B1(new_n434), .B2(new_n386), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n669), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n403), .A2(new_n418), .ZN(new_n878));
  INV_X1    g0678(.A(new_n669), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n403), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n437), .ZN(new_n882));
  INV_X1    g0682(.A(new_n437), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n421), .B2(new_n669), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n876), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n886), .C1(new_n442), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n873), .B(KEYINPUT39), .C1(new_n887), .C2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n437), .B1(new_n420), .B2(new_n421), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n420), .A2(new_n669), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n882), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT106), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n895), .A2(new_n898), .A3(new_n882), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n419), .A2(new_n439), .A3(new_n422), .A4(new_n440), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n894), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n892), .B(new_n889), .C1(new_n902), .C2(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n891), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n886), .B1(new_n442), .B2(new_n888), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n892), .B1(new_n907), .B2(new_n889), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n873), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n872), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n832), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n704), .B2(new_n834), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n316), .A2(new_n671), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n343), .A2(new_n348), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n329), .A2(new_n332), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(new_n339), .A3(new_n341), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n316), .B(new_n671), .C1(new_n916), .C2(new_n347), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n907), .A2(new_n889), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n423), .B2(new_n669), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT92), .B1(new_n719), .B2(new_n672), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n709), .B(new_n671), .C1(new_n718), .C2(new_n655), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT29), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT93), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n721), .A2(new_n708), .A3(KEYINPUT29), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n706), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n443), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n638), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n923), .B(new_n931), .Z(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n887), .A2(new_n890), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n833), .B1(new_n914), .B2(new_n917), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n742), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n742), .A2(KEYINPUT40), .A3(new_n935), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n896), .A2(KEYINPUT106), .B1(new_n894), .B2(new_n900), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n940), .B2(new_n899), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n941), .B2(new_n890), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n930), .A2(new_n742), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(G330), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n932), .A2(KEYINPUT107), .A3(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(new_n209), .B2(new_n747), .C1(new_n932), .C2(new_n947), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT107), .B1(new_n932), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n871), .B1(new_n949), .B2(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n611), .A2(new_n671), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n618), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n658), .B2(new_n952), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT108), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n544), .B1(new_n535), .B2(new_n672), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n650), .A2(new_n671), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n692), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n543), .B1(new_n958), .B2(new_n628), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n962), .A2(KEYINPUT42), .B1(new_n672), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n957), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n955), .A2(new_n956), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n687), .A2(new_n961), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n695), .B(KEYINPUT41), .Z(new_n971));
  INV_X1    g0771(.A(new_n691), .ZN(new_n972));
  INV_X1    g0772(.A(new_n686), .ZN(new_n973));
  INV_X1    g0773(.A(new_n681), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n692), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n676), .A2(KEYINPUT110), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n725), .A2(new_n743), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n692), .A2(new_n684), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n960), .B1(KEYINPUT109), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT109), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n981), .A2(new_n987), .A3(new_n983), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n692), .A2(new_n684), .A3(new_n960), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n687), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AND4_X1   g0793(.A1(new_n687), .A2(new_n992), .A3(new_n986), .A4(new_n988), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT111), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n725), .A2(new_n996), .A3(new_n743), .A4(new_n978), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n980), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n971), .B1(new_n998), .B2(new_n744), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n970), .B1(new_n999), .B2(new_n749), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n823), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n955), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n256), .B1(new_n771), .B2(G317), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n796), .B2(new_n456), .ZN(new_n1004));
  INV_X1    g0804(.A(G283), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n789), .A2(new_n1005), .B1(new_n790), .B2(new_n205), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G107), .C2(new_n778), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT46), .B1(new_n782), .B2(G116), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n782), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G311), .C2(new_n765), .ZN(new_n1010));
  INV_X1    g0810(.A(G294), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1007), .B(new_n1010), .C1(new_n1011), .C2(new_n804), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n778), .A2(G68), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n796), .B2(new_n275), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n765), .A2(G143), .B1(new_n1014), .B2(KEYINPUT112), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(KEYINPUT112), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n789), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(G50), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n252), .B1(new_n771), .B2(G137), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n781), .A2(G77), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n782), .A2(G58), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n804), .B2(new_n798), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT47), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n807), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n816), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n814), .B1(new_n213), .B2(new_n355), .C1(new_n1028), .C2(new_n238), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1002), .A2(new_n750), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1000), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n980), .A2(new_n997), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n695), .C1(new_n744), .C2(new_n978), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n978), .A2(new_n749), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT113), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1001), .B1(new_n973), .B2(new_n974), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n350), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT50), .B1(new_n350), .B2(new_n202), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n697), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n816), .B(new_n1040), .C1(new_n235), .C2(new_n446), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n819), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(G107), .B2(new_n213), .C1(new_n697), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n751), .B1(new_n1043), .B2(new_n814), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT114), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n252), .B1(new_n785), .B2(G68), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n275), .B2(new_n770), .C1(new_n796), .C2(new_n202), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n255), .A2(new_n792), .B1(new_n790), .B2(new_n205), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n354), .C2(new_n778), .ZN(new_n1049));
  INV_X1    g0849(.A(G159), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n764), .C1(new_n273), .C2(new_n804), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n256), .B1(new_n771), .B2(G326), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1017), .A2(G303), .B1(G317), .B2(new_n767), .ZN(new_n1053));
  INV_X1    g0853(.A(G322), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n764), .C1(new_n804), .C2(new_n773), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n782), .A2(G294), .B1(G283), .B2(new_n778), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT115), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1052), .B1(new_n466), .B2(new_n790), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1051), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1045), .B1(new_n1065), .B2(new_n807), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1035), .B1(new_n1036), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1033), .A2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n995), .A2(new_n749), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n814), .B1(new_n205), .B2(new_n213), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n243), .B2(new_n816), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n252), .B1(new_n770), .B2(new_n1054), .C1(new_n1011), .C2(new_n774), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G116), .B2(new_n778), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G107), .A2(new_n781), .B1(new_n782), .B2(G283), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n804), .C2(new_n456), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n765), .A2(G317), .B1(G311), .B2(new_n767), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n761), .A2(G50), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n778), .A2(G77), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n252), .B1(new_n771), .B2(G143), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n847), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1017), .A2(new_n350), .B1(G68), .B2(new_n782), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n764), .A2(new_n275), .B1(new_n1050), .B2(new_n796), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n1075), .A2(new_n1077), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n751), .B(new_n1071), .C1(new_n1086), .C2(new_n807), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n813), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n960), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n998), .A2(new_n695), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n995), .B1(new_n980), .B2(new_n997), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1069), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(G390));
  OR2_X1    g0892(.A1(new_n908), .A2(new_n873), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n872), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n912), .B2(new_n919), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1093), .A2(new_n1095), .A3(new_n903), .A4(new_n891), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n831), .B(new_n918), .C1(new_n721), .C2(new_n911), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n889), .B1(new_n902), .B2(KEYINPUT38), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n742), .A2(G330), .A3(new_n834), .A4(new_n918), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n748), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n750), .B1(new_n350), .B2(new_n856), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n904), .A2(new_n909), .A3(new_n812), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n793), .A2(new_n256), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT117), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n789), .A2(new_n205), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n771), .A2(G294), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n767), .A2(G116), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n838), .A2(new_n1079), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1108), .B(new_n1111), .C1(G283), .C2(new_n765), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1107), .B(new_n1112), .C1(new_n206), .C2(new_n804), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT118), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n804), .A2(new_n842), .ZN(new_n1116));
  INV_X1    g0916(.A(G125), .ZN(new_n1117));
  INV_X1    g0917(.A(G132), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n256), .B1(new_n770), .B2(new_n1117), .C1(new_n796), .C2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n789), .A2(new_n1120), .B1(new_n790), .B2(new_n202), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G159), .C2(new_n778), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n782), .A2(G150), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT53), .Z(new_n1124));
  NAND2_X1  g0924(.A1(new_n765), .A2(G128), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n1116), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1104), .B(new_n1105), .C1(new_n807), .C2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1103), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT116), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n443), .A2(new_n743), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n742), .A2(G330), .A3(new_n834), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n919), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1100), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n663), .A2(new_n672), .A3(new_n834), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n832), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n831), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n924), .A2(new_n925), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n832), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n1136), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n931), .A2(new_n1132), .A3(new_n1133), .A4(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n930), .B(new_n707), .C1(new_n722), .C2(new_n724), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(new_n1143), .A3(new_n639), .A4(new_n1133), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1100), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n872), .B1(new_n1138), .B2(new_n918), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1152), .A2(new_n904), .A3(new_n909), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1099), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AND4_X1   g0955(.A1(new_n639), .A2(new_n1145), .A3(new_n1143), .A4(new_n1133), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n695), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1131), .B1(new_n1150), .B2(new_n1159), .ZN(G378));
  AOI21_X1  g0960(.A(new_n936), .B1(new_n907), .B2(new_n889), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n942), .B(G330), .C1(new_n1161), .C2(KEYINPUT40), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n294), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n305), .A2(new_n1163), .A3(new_n879), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n293), .B1(new_n294), .B2(new_n669), .C1(new_n303), .C2(new_n304), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(KEYINPUT121), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n937), .A2(G330), .A3(new_n942), .A4(new_n1171), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n923), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n910), .A3(new_n1174), .A4(new_n922), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT122), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(KEYINPUT122), .A3(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1169), .A2(new_n811), .A3(new_n1170), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G58), .A2(new_n781), .B1(new_n782), .B2(G77), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n252), .A2(new_n264), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n767), .B2(G107), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n354), .A2(new_n785), .B1(new_n771), .B2(G283), .ZN(new_n1187));
  AND4_X1   g0987(.A1(new_n1013), .A2(new_n1184), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n466), .B2(new_n764), .C1(new_n804), .C2(new_n205), .ZN(new_n1189));
  XOR2_X1   g0989(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1190));
  OR2_X1    g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1185), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G128), .A2(new_n767), .B1(new_n778), .B2(G150), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n792), .B2(new_n1120), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n761), .A2(G132), .B1(G137), .B2(new_n785), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT120), .Z(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G125), .C2(new_n765), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n771), .C2(G124), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n790), .B2(new_n798), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(KEYINPUT59), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1194), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n807), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n750), .B1(G50), .B2(new_n856), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1182), .A2(new_n748), .B1(new_n1183), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n931), .A2(new_n1133), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1182), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1178), .A2(KEYINPUT57), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1158), .A2(new_n931), .A3(new_n1133), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n696), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1208), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(G375));
  NAND2_X1  g1018(.A1(new_n919), .A2(new_n811), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n750), .B1(G68), .B2(new_n856), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT123), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n767), .A2(G137), .B1(G128), .B2(new_n771), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n256), .C1(new_n275), .C2(new_n774), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n380), .A2(new_n790), .B1(new_n792), .B2(new_n1050), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G50), .C2(new_n778), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n1118), .B2(new_n764), .C1(new_n804), .C2(new_n1120), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n796), .A2(new_n1005), .B1(new_n355), .B2(new_n777), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1227), .A2(new_n1228), .B1(new_n1011), .B2(new_n764), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1228), .B2(new_n1227), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n789), .A2(new_n206), .B1(new_n792), .B2(new_n205), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1020), .B(new_n252), .C1(new_n456), .C2(new_n770), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1230), .B(new_n1233), .C1(new_n466), .C2(new_n804), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1226), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1221), .B1(new_n1235), .B2(new_n807), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1143), .A2(new_n749), .B1(new_n1219), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1143), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1210), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n971), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1237), .B1(new_n1241), .B2(new_n1148), .ZN(G381));
  NAND3_X1  g1042(.A1(new_n1033), .A2(new_n827), .A3(new_n1067), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(G384), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1244), .A2(G390), .A3(G378), .A4(G381), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1245), .A2(new_n1000), .A3(new_n1030), .A4(new_n1217), .ZN(G407));
  INV_X1    g1046(.A(G378), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1217), .A2(new_n670), .A3(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(G213), .A3(new_n1248), .ZN(G409));
  AND3_X1   g1049(.A1(new_n1000), .A2(new_n1030), .A3(G390), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G390), .B1(new_n1000), .B2(new_n1030), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT127), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1243), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(KEYINPUT127), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1207), .A2(new_n1183), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1176), .A2(KEYINPUT122), .A3(new_n1177), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT122), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1260), .B1(new_n1263), .B2(new_n749), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1263), .B2(new_n1215), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n695), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1264), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1215), .A2(new_n1240), .A3(new_n1181), .A4(new_n1180), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1260), .B1(new_n1178), .B2(new_n749), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1247), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1146), .A2(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1239), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1210), .A2(KEYINPUT60), .A3(new_n1238), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n695), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G384), .A3(new_n1237), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1276), .B2(new_n1237), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(G343), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1272), .A2(new_n1280), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1272), .A2(KEYINPUT125), .A3(new_n1280), .A4(new_n1283), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT62), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1272), .A2(new_n1283), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1279), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(G2897), .A3(new_n1277), .A4(new_n1282), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1282), .A2(G2897), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1259), .B1(new_n1288), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1280), .A4(new_n1283), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1258), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT63), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1286), .A2(new_n1302), .A3(new_n1287), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1289), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1283), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1294), .A3(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1301), .A2(new_n1303), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1298), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1247), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1258), .A2(new_n1267), .A3(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1217), .B(G378), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n1257), .A3(new_n1255), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1311), .A2(new_n1280), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1280), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(G402));
endmodule


