//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  OR2_X1    g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n193), .A3(new_n188), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n200), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(G134), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n203), .ZN(new_n208));
  AOI211_X1 g022(.A(G131), .B(new_n202), .C1(new_n205), .C2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n208), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n199), .A2(new_n201), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n197), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G119), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n220), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n215), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n207), .B1(new_n206), .B2(new_n203), .ZN(new_n227));
  AOI211_X1 g041(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n198), .C2(G134), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n212), .B(new_n210), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n194), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n191), .A2(new_n193), .A3(new_n233), .A4(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n206), .A2(new_n201), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n214), .A2(new_n226), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n214), .A2(new_n241), .A3(new_n226), .A4(new_n238), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT31), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n191), .A2(new_n193), .B1(new_n187), .B2(new_n188), .ZN(new_n247));
  INV_X1    g061(.A(new_n196), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n212), .B1(new_n227), .B2(new_n228), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G131), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n249), .B1(new_n251), .B2(new_n229), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n229), .A2(new_n235), .A3(new_n237), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n246), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n214), .A2(KEYINPUT30), .A3(new_n238), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n225), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n257), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n243), .A2(new_n244), .A3(new_n256), .A4(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n256), .A2(new_n240), .A3(new_n242), .A4(new_n263), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT31), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n239), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n225), .B1(new_n252), .B2(new_n253), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n240), .A2(new_n242), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n271), .B2(KEYINPUT28), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n264), .B(new_n266), .C1(new_n272), .C2(new_n263), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n274));
  NOR2_X1   g088(.A1(G472), .A2(G902), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(KEYINPUT28), .ZN(new_n278));
  INV_X1    g092(.A(new_n263), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n268), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n243), .A2(new_n256), .A3(new_n279), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n272), .B2(new_n279), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G472), .ZN(new_n288));
  OAI22_X1  g102(.A1(new_n276), .A2(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n273), .A2(new_n275), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n286), .A2(new_n280), .ZN(new_n296));
  OAI21_X1  g110(.A(G472), .B1(new_n296), .B2(new_n284), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(KEYINPUT68), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n217), .A2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT24), .B(G110), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT23), .B1(new_n299), .B2(G119), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(KEYINPUT69), .A3(KEYINPUT23), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n299), .A3(G119), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT70), .B1(new_n217), .B2(G128), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n307), .A2(new_n308), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(new_n300), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n304), .B1(new_n314), .B2(G110), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G140), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT72), .A2(G125), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT72), .A2(G125), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n321), .B2(G140), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NOR4_X1   g137(.A1(new_n319), .A2(new_n320), .A3(new_n316), .A4(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT16), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT16), .A2(G140), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n319), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n329), .B(new_n326), .C1(new_n319), .C2(new_n320), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(G146), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n190), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n315), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n302), .A2(new_n303), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g151(.A(new_n318), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT72), .B(G125), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n323), .ZN(new_n340));
  OR2_X1    g154(.A1(KEYINPUT72), .A2(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT72), .A2(G125), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(KEYINPUT73), .A3(G140), .A4(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n337), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n329), .B1(new_n339), .B2(new_n326), .ZN(new_n345));
  INV_X1    g159(.A(new_n330), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n190), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n336), .B1(new_n348), .B2(new_n332), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n300), .A2(new_n313), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n311), .A2(new_n310), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT69), .B1(new_n301), .B2(KEYINPUT23), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n351), .B1(new_n354), .B2(new_n308), .ZN(new_n355));
  INV_X1    g169(.A(G110), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT71), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n314), .A2(new_n358), .A3(G110), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n349), .A2(new_n350), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n350), .B1(new_n349), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n335), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT76), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT22), .B(G137), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n335), .B(new_n367), .C1(new_n361), .C2(new_n362), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G234), .B2(new_n283), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n283), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n371), .A2(KEYINPUT25), .A3(new_n283), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n376), .B1(new_n381), .B2(new_n373), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n291), .A2(new_n298), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G210), .B1(G237), .B2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n235), .A2(new_n321), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n259), .A2(G224), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n197), .A2(new_n339), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n339), .B1(new_n232), .B2(new_n234), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n321), .B1(new_n195), .B2(new_n196), .ZN(new_n393));
  OAI211_X1 g207(.A(G224), .B(new_n259), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n217), .A3(G116), .ZN(new_n399));
  OAI211_X1 g213(.A(G113), .B(new_n399), .C1(new_n223), .C2(new_n398), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n222), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT3), .B1(new_n402), .B2(G107), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  INV_X1    g218(.A(G107), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(G104), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(G107), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n402), .A2(G107), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n405), .A2(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n409), .A2(new_n412), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n222), .A3(new_n400), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT8), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n388), .A2(new_n390), .A3(new_n395), .A4(new_n389), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n397), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G101), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT4), .A3(new_n409), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(G101), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n225), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n418), .A3(new_n416), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n422), .ZN(new_n432));
  INV_X1    g246(.A(new_n419), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n414), .B2(new_n416), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n421), .B1(new_n435), .B2(new_n397), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n283), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n416), .ZN(new_n438));
  INV_X1    g252(.A(new_n418), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n391), .A2(new_n394), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n443), .A3(new_n439), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n387), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n397), .A2(new_n420), .A3(new_n422), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n430), .A3(new_n423), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(new_n283), .A3(new_n386), .A4(new_n445), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n385), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n453));
  NOR2_X1   g267(.A1(G475), .A2(G902), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n455));
  OAI211_X1 g269(.A(G146), .B(new_n343), .C1(new_n455), .C2(new_n318), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n334), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT83), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n459), .A3(new_n334), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n258), .A2(new_n259), .A3(G214), .ZN(new_n461));
  NOR2_X1   g275(.A1(KEYINPUT82), .A2(G143), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(KEYINPUT82), .A2(G143), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n461), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n458), .A2(new_n460), .A3(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT19), .B(new_n343), .C1(new_n455), .C2(new_n318), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT19), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n333), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n190), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n463), .A2(G131), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n467), .A2(new_n210), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n332), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n190), .A3(new_n475), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n471), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n402), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(KEYINPUT85), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n477), .A2(new_n478), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n463), .A2(KEYINPUT17), .A3(G131), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n348), .A2(new_n489), .A3(new_n332), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n485), .A3(new_n471), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT85), .B1(new_n483), .B2(new_n486), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n454), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT20), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(new_n454), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT86), .B(G475), .Z(new_n500));
  AOI21_X1  g314(.A(new_n485), .B1(new_n491), .B2(new_n471), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n492), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n501), .B2(KEYINPUT87), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G478), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n192), .A2(G128), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n299), .A2(G143), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G134), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n200), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G116), .B(G122), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n405), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n219), .A2(KEYINPUT14), .A3(G122), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(G107), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(KEYINPUT88), .A3(G107), .A4(new_n520), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n515), .B(new_n405), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n509), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n510), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n509), .A2(new_n527), .ZN(new_n530));
  OAI21_X1  g344(.A(G134), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n531), .A3(new_n513), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT9), .B(G234), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n534), .A2(new_n372), .A3(G953), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OR3_X1    g350(.A1(new_n525), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n525), .B2(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT15), .B(new_n508), .C1(new_n539), .C2(new_n283), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n541));
  AOI211_X1 g355(.A(G902), .B(new_n541), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  INV_X1    g356(.A(G952), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G953), .ZN(new_n544));
  NAND2_X1  g358(.A1(G234), .A2(G237), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n545), .A2(G902), .A3(G953), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT21), .B(G898), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n540), .A2(new_n542), .A3(new_n549), .ZN(new_n550));
  AND4_X1   g364(.A1(new_n453), .A2(new_n499), .A3(new_n507), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n506), .B1(new_n496), .B2(new_n498), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n453), .B1(new_n552), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n452), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n555));
  INV_X1    g369(.A(new_n234), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n191), .A2(new_n558), .A3(KEYINPUT1), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(G128), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n556), .B1(new_n560), .B2(new_n194), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n555), .B1(new_n561), .B2(new_n413), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n209), .A2(new_n213), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n426), .A2(new_n197), .A3(new_n428), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n415), .A2(new_n235), .A3(KEYINPUT10), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n413), .A2(new_n232), .A3(new_n234), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n561), .B2(new_n413), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n251), .A2(new_n229), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n568), .A2(KEYINPUT12), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT12), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(G110), .B(G140), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT77), .ZN(new_n574));
  INV_X1    g388(.A(G227), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n574), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n569), .ZN(new_n580));
  INV_X1    g394(.A(new_n577), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n566), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G469), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT79), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n581), .A2(new_n566), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n572), .A2(new_n577), .B1(new_n587), .B2(new_n580), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n586), .B(G469), .C1(new_n588), .C2(G902), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n570), .A2(new_n571), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n590), .A2(new_n587), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n581), .B1(new_n580), .B2(new_n566), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n584), .B(new_n283), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n585), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT80), .ZN(new_n595));
  OAI21_X1  g409(.A(G221), .B1(new_n534), .B2(G902), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n554), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n383), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  AOI21_X1  g416(.A(KEYINPUT25), .B1(new_n371), .B2(new_n283), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n378), .B(G902), .C1(new_n369), .C2(new_n370), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n373), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n264), .A2(new_n266), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n263), .B1(new_n278), .B2(new_n268), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n283), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n608), .A2(G472), .B1(new_n275), .B2(new_n273), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n549), .B(new_n385), .C1(new_n447), .C2(new_n451), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n375), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n599), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(G478), .B1(new_n539), .B2(new_n283), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT90), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(KEYINPUT90), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n539), .B(KEYINPUT33), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n508), .A2(G902), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n614), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n552), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  XNOR2_X1  g436(.A(new_n499), .B(KEYINPUT91), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n507), .B1(new_n540), .B2(new_n542), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n612), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NAND2_X1  g443(.A1(new_n447), .A2(new_n451), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n384), .ZN(new_n631));
  INV_X1    g445(.A(new_n498), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n483), .A2(new_n486), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT85), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n492), .A3(new_n487), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n497), .B1(new_n636), .B2(new_n454), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n550), .B(new_n507), .C1(new_n632), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT89), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n552), .A2(new_n453), .A3(new_n550), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n594), .A2(new_n596), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT80), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n265), .B(new_n244), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n278), .A2(new_n268), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n279), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n292), .B1(new_n649), .B2(new_n288), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n363), .A2(KEYINPUT92), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n363), .A2(KEYINPUT92), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n363), .A2(KEYINPUT92), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n374), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n650), .B1(new_n605), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n641), .A2(new_n645), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n605), .A2(new_n659), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n645), .A2(new_n291), .A3(new_n298), .A4(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n546), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n547), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n665), .A2(new_n625), .A3(new_n631), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n299), .ZN(G30));
  INV_X1    g486(.A(new_n664), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n630), .B(KEYINPUT38), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n384), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n540), .A2(new_n542), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n552), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n279), .B1(new_n243), .B2(new_n256), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n283), .B1(new_n271), .B2(new_n263), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n295), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n675), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT93), .B(KEYINPUT39), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n669), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n645), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NAND2_X1  g504(.A1(new_n619), .A2(new_n669), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT94), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT94), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n619), .A2(new_n693), .A3(new_n669), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n665), .A2(new_n695), .A3(new_n631), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT95), .B(G146), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G48));
  NAND2_X1  g512(.A1(new_n580), .A2(new_n566), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n590), .A2(new_n587), .B1(new_n699), .B2(new_n577), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n593), .A2(new_n701), .A3(new_n596), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n291), .A2(new_n298), .A3(new_n382), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n619), .A3(new_n610), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT41), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G113), .ZN(G15));
  NAND3_X1  g521(.A1(new_n704), .A2(new_n610), .A3(new_n626), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND3_X1  g523(.A1(new_n291), .A2(new_n298), .A3(new_n664), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n639), .A2(new_n640), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n631), .A2(KEYINPUT96), .A3(new_n702), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT96), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n703), .B2(new_n452), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n711), .A2(KEYINPUT97), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT97), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n712), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(new_n710), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT98), .B(G119), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G21));
  INV_X1    g537(.A(KEYINPUT100), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n647), .A2(KEYINPUT99), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT99), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n279), .B1(new_n272), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n646), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n728), .A2(new_n275), .B1(new_n608), .B2(G472), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n382), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n605), .A2(new_n375), .ZN(new_n731));
  INV_X1    g545(.A(new_n729), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT100), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NOR4_X1   g548(.A1(new_n677), .A2(new_n549), .A3(new_n631), .A4(new_n702), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NAND2_X1  g551(.A1(new_n664), .A2(new_n729), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT101), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n664), .A2(KEYINPUT101), .A3(new_n729), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n695), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n716), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  INV_X1    g559(.A(new_n593), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n583), .A2(new_n584), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n596), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n385), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n447), .A2(new_n451), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n291), .A2(new_n298), .A3(new_n382), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n695), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n731), .B1(new_n297), .B2(new_n295), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT42), .A3(new_n752), .ZN(new_n756));
  OAI22_X1  g570(.A1(new_n754), .A2(KEYINPUT42), .B1(new_n756), .B2(new_n695), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT102), .B(G131), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G33));
  NOR2_X1   g573(.A1(new_n625), .A2(new_n670), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n383), .A3(new_n752), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n578), .A2(new_n582), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT104), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n584), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT103), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT105), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n746), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n749), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n685), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n630), .A2(new_n385), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n552), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  OAI22_X1  g597(.A1(new_n782), .A2(new_n618), .B1(KEYINPUT106), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n618), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n552), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n650), .A3(new_n664), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n198), .ZN(G39));
  OR2_X1    g608(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n781), .B(new_n382), .C1(new_n291), .C2(new_n298), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n743), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  AND2_X1   g614(.A1(new_n788), .A2(new_n546), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n593), .A2(new_n701), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n751), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n755), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT48), .Z(new_n807));
  AND2_X1   g621(.A1(new_n801), .A2(new_n734), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n716), .ZN(new_n809));
  INV_X1    g623(.A(new_n619), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n682), .A2(new_n382), .A3(new_n546), .A4(new_n803), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n809), .B(new_n544), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n807), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n674), .A2(new_n384), .A3(new_n702), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT50), .Z(new_n819));
  NOR3_X1   g633(.A1(new_n811), .A2(new_n782), .A3(new_n785), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n805), .B2(new_n742), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n808), .A2(new_n780), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n795), .A2(new_n796), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n593), .A2(new_n701), .A3(new_n749), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n816), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n827), .B(KEYINPUT118), .Z(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n832), .B2(new_n822), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT120), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n828), .A2(new_n830), .A3(new_n822), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n833), .A4(new_n816), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n641), .A2(new_n645), .A3(new_n660), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n552), .B1(new_n540), .B2(new_n542), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n599), .A2(new_n611), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT109), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n383), .A2(new_n600), .B1(new_n612), .B2(new_n619), .ZN(new_n845));
  INV_X1    g659(.A(new_n611), .ZN(new_n846));
  INV_X1    g660(.A(new_n842), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n645), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT109), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n661), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT110), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT108), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n717), .A2(new_n720), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n708), .A2(new_n705), .A3(new_n736), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n705), .A2(new_n736), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(KEYINPUT108), .A3(new_n721), .A4(new_n708), .ZN(new_n861));
  INV_X1    g675(.A(new_n665), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n507), .A2(new_n676), .A3(new_n669), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n623), .A2(new_n781), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n692), .A2(new_n694), .A3(new_n752), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n862), .A2(new_n864), .B1(new_n742), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n757), .A2(new_n866), .A3(new_n761), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n855), .A2(new_n859), .A3(new_n861), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n665), .A2(new_n631), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n760), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n743), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n677), .A2(new_n631), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n681), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n669), .A2(KEYINPUT112), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n669), .A2(KEYINPUT112), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n749), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n746), .B2(new_n747), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n664), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT113), .B1(new_n664), .B2(new_n877), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n870), .A2(new_n871), .A3(new_n881), .A4(new_n744), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n716), .A2(new_n692), .A3(new_n694), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n741), .B2(new_n740), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n671), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n696), .A2(new_n880), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT52), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n840), .B1(new_n868), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n857), .A2(new_n858), .A3(new_n840), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n855), .A2(new_n894), .A3(new_n867), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT111), .B1(new_n671), .B2(new_n886), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT111), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n870), .A2(new_n897), .A3(new_n744), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n880), .A2(new_n883), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n896), .A2(new_n898), .A3(new_n871), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n882), .A2(new_n883), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT114), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT114), .B1(new_n900), .B2(new_n901), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  OAI211_X1 g721(.A(KEYINPUT117), .B(new_n840), .C1(new_n868), .C2(new_n890), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n893), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n868), .ZN(new_n910));
  INV_X1    g724(.A(new_n890), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(KEYINPUT53), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT115), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n910), .A2(new_n914), .A3(new_n911), .A4(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n902), .B(new_n903), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT53), .B1(new_n917), .B2(new_n910), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT116), .B(new_n909), .C1(new_n919), .C2(new_n907), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(KEYINPUT54), .C1(new_n916), .C2(new_n918), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n839), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n382), .A2(new_n750), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT107), .Z(new_n926));
  XNOR2_X1  g740(.A(new_n802), .B(KEYINPUT49), .ZN(new_n927));
  OR4_X1    g741(.A1(new_n674), .A2(new_n681), .A3(new_n786), .A4(new_n927), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n923), .A2(new_n924), .B1(new_n926), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n259), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n893), .A2(new_n908), .A3(new_n906), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n441), .A2(new_n444), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n442), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT56), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n940), .B2(new_n933), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n942), .B2(new_n937), .ZN(G51));
  INV_X1    g757(.A(new_n932), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n944), .A2(new_n283), .A3(new_n771), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n909), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n772), .B(KEYINPUT122), .Z(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT57), .Z(new_n949));
  AOI21_X1  g763(.A(new_n700), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n949), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n946), .B2(new_n909), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT123), .B1(new_n954), .B2(new_n700), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n930), .B1(new_n952), .B2(new_n955), .ZN(G54));
  NOR2_X1   g770(.A1(new_n944), .A2(new_n283), .ZN(new_n957));
  AND2_X1   g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n957), .A2(new_n636), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n636), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n930), .ZN(G60));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n947), .A2(new_n616), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n931), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n920), .A2(new_n922), .A3(new_n964), .ZN(new_n967));
  INV_X1    g781(.A(new_n616), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n370), .B(new_n369), .C1(new_n944), .C2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n932), .B(new_n973), .C1(new_n656), .C2(new_n658), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n931), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  INV_X1    g791(.A(new_n548), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n259), .B1(new_n978), .B2(G224), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n855), .A2(new_n859), .A3(new_n861), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n259), .ZN(new_n981));
  INV_X1    g795(.A(G898), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n935), .B1(new_n982), .B2(G953), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n981), .B(new_n983), .ZN(G69));
  NAND2_X1  g798(.A1(new_n472), .A2(new_n475), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT124), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n254), .A2(new_n255), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  NAND2_X1  g803(.A1(G900), .A2(G953), .ZN(new_n990));
  INV_X1    g804(.A(new_n779), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n755), .A2(new_n872), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n793), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n757), .A2(new_n761), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n896), .A2(new_n871), .A3(new_n898), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n799), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n989), .B(new_n990), .C1(new_n996), .C2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n689), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n781), .B1(new_n810), .B2(new_n842), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n383), .A2(new_n645), .A3(new_n685), .A4(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n793), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n999), .A2(new_n799), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1004), .A2(new_n259), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n997), .B1(new_n1005), .B2(new_n989), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n575), .B2(new_n667), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n989), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1006), .B(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n1004), .B2(new_n980), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1015), .A2(new_n678), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n285), .A2(new_n1012), .ZN(new_n1018));
  OR3_X1    g832(.A1(new_n919), .A2(new_n678), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1012), .B1(new_n996), .B2(new_n980), .ZN(new_n1020));
  INV_X1    g834(.A(new_n285), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n930), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1017), .A2(new_n1019), .A3(new_n1022), .ZN(G57));
endmodule


