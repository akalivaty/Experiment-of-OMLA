//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G50), .A2(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n203), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI211_X1 g0016(.A(new_n214), .B(new_n216), .C1(G77), .C2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n204), .A2(new_n205), .ZN(new_n231));
  INV_X1    g0031(.A(G50), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n211), .B(new_n227), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G226), .B(G232), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n221), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n202), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n228), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT11), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n229), .A2(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G13), .ZN(new_n268));
  OR3_X1    g0068(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT12), .B1(new_n268), .B2(G68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n252), .A2(new_n267), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(G68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G226), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G97), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(G232), .A4(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n278), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n276), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G238), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(new_n291), .B2(new_n295), .ZN(new_n297));
  OAI21_X1  g0097(.A(G200), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G190), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n274), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n296), .A2(new_n297), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n306), .B2(G179), .ZN(new_n310));
  OAI211_X1 g0110(.A(G169), .B(new_n304), .C1(new_n296), .C2(new_n297), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n303), .B1(new_n312), .B2(new_n273), .ZN(new_n313));
  INV_X1    g0113(.A(G244), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n293), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n278), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n283), .A2(new_n285), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT67), .B1(new_n318), .B2(new_n280), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT67), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n279), .A2(new_n320), .A3(G1698), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n213), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n279), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G232), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n318), .A2(new_n325), .A3(G1698), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n316), .B(new_n317), .C1(new_n327), .C2(new_n289), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(G179), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n268), .A2(G77), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n271), .A2(G77), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n229), .A2(new_n260), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n333), .A2(new_n334), .B1(new_n229), .B2(new_n263), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n336), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n262), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n252), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n331), .B(new_n332), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n328), .A2(new_n307), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n329), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n317), .B1(new_n327), .B2(new_n289), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  OR3_X1    g0147(.A1(new_n346), .A2(new_n347), .A3(new_n315), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n328), .B2(G200), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n352));
  INV_X1    g0152(.A(G150), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n333), .A2(new_n262), .B1(new_n353), .B2(new_n334), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n257), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G13), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n356), .A2(new_n229), .A3(G1), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n232), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n267), .B1(new_n254), .B2(new_n255), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G50), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n355), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n361), .A2(KEYINPUT9), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(KEYINPUT9), .ZN(new_n363));
  INV_X1    g0163(.A(G223), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n319), .B2(new_n321), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n279), .A2(G222), .A3(new_n280), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n263), .B2(new_n279), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n290), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n294), .A2(G226), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n317), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n362), .A2(new_n363), .B1(G200), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(new_n347), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n370), .B2(G200), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n362), .A2(new_n363), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(G200), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n372), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n375), .A2(new_n373), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n370), .A2(new_n307), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n361), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT69), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT69), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n386), .A3(new_n361), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n385), .B(new_n387), .C1(G179), .C2(new_n370), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n313), .A2(new_n351), .A3(new_n382), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT77), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n268), .A2(new_n333), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n359), .B2(new_n333), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT76), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n318), .B2(new_n229), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n396), .B(G20), .C1(new_n283), .C2(new_n285), .ZN(new_n397));
  OAI21_X1  g0197(.A(G68), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n204), .A2(new_n205), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT73), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n334), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n258), .A2(KEYINPUT73), .A3(G159), .ZN(new_n404));
  AOI22_X1  g0204(.A1(G20), .A2(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT74), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n398), .A2(KEYINPUT74), .A3(KEYINPUT16), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n284), .A2(KEYINPUT75), .A3(G33), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n283), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT75), .B1(new_n284), .B2(G33), .ZN(new_n413));
  OAI211_X1 g0213(.A(KEYINPUT7), .B(new_n229), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n396), .B1(new_n279), .B2(G20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G68), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n405), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n342), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n394), .B1(new_n410), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n364), .A2(new_n280), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n279), .B(new_n422), .C1(G226), .C2(new_n280), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n289), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n317), .B1(new_n293), .B2(new_n325), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G179), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n307), .B2(new_n427), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n391), .B1(new_n421), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n203), .B1(new_n414), .B2(new_n415), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n400), .A2(G20), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n403), .A2(new_n404), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n419), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n252), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n408), .B2(new_n409), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT18), .B(new_n429), .C1(new_n438), .C2(new_n394), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n284), .A2(G33), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n442));
  OAI211_X1 g0242(.A(KEYINPUT7), .B(new_n229), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n203), .B1(new_n415), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n435), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT74), .B1(new_n445), .B2(KEYINPUT16), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n444), .A2(new_n435), .A3(new_n407), .A4(new_n419), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n252), .B(new_n436), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(G200), .B1(new_n425), .B2(new_n426), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n427), .A2(G190), .ZN(new_n450));
  INV_X1    g0250(.A(new_n394), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n449), .A4(new_n450), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n390), .B1(new_n440), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n456), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n431), .A2(new_n439), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n389), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n219), .A2(new_n280), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n224), .A2(G1698), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n283), .A2(new_n462), .A3(new_n285), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G294), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n290), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(G41), .ZN(new_n470));
  INV_X1    g0270(.A(G41), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n470), .A2(new_n472), .A3(new_n474), .A4(G274), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(new_n474), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G264), .A3(new_n289), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n467), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G169), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT89), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n467), .A2(G179), .A3(new_n475), .A4(new_n477), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n479), .B2(new_n481), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n283), .A2(new_n285), .A3(new_n229), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n279), .A2(new_n229), .A3(G87), .A4(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n229), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT23), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT82), .B(G116), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n261), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n488), .A2(new_n489), .B1(new_n494), .B2(new_n261), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n492), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n342), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT88), .B1(new_n268), .B2(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT88), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n357), .A2(new_n503), .A3(new_n323), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT25), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n267), .A2(G13), .B1(new_n275), .B2(G33), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n256), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n323), .B2(new_n511), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n483), .A2(new_n484), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n501), .A2(new_n512), .ZN(new_n514));
  INV_X1    g0314(.A(G200), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n478), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G190), .B2(new_n478), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n219), .B1(new_n473), .B2(G1), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n275), .A2(new_n277), .A3(G45), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n289), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n213), .A2(new_n280), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n314), .A2(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n283), .A2(new_n524), .A3(new_n285), .A4(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(KEYINPUT82), .A2(G116), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT82), .A2(G116), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(G33), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n523), .B1(new_n531), .B2(new_n290), .ZN(new_n532));
  INV_X1    g0332(.A(G179), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n289), .B1(new_n526), .B2(new_n530), .ZN(new_n535));
  NOR4_X1   g0335(.A1(new_n535), .A2(new_n523), .A3(KEYINPUT83), .A4(G179), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n535), .A2(new_n523), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n307), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n339), .A2(new_n357), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n218), .A2(new_n223), .A3(new_n323), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n282), .A2(new_n229), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT19), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n283), .A2(new_n285), .A3(new_n229), .A4(G68), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n282), .B2(G20), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n252), .ZN(new_n549));
  XOR2_X1   g0349(.A(new_n339), .B(KEYINPUT84), .Z(new_n550));
  OAI211_X1 g0350(.A(new_n541), .B(new_n549), .C1(new_n550), .C2(new_n511), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n540), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n532), .A2(G190), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n515), .B2(new_n532), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n256), .A2(G87), .A3(new_n510), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n549), .A2(new_n556), .A3(new_n541), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n538), .A2(new_n552), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n513), .A2(new_n518), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT86), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT20), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n493), .A2(G20), .B1(new_n228), .B2(new_n251), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n567), .B(new_n229), .C1(G33), .C2(new_n223), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(KEYINPUT82), .A2(G116), .ZN(new_n570));
  OAI21_X1  g0370(.A(G20), .B1(new_n570), .B2(new_n527), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n252), .A3(new_n568), .ZN(new_n572));
  INV_X1    g0372(.A(new_n565), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n564), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n493), .A2(new_n357), .ZN(new_n576));
  INV_X1    g0376(.A(new_n510), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n577), .A2(new_n220), .A3(new_n252), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G264), .A2(G1698), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n279), .B(new_n581), .C1(new_n224), .C2(G1698), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n289), .B1(new_n318), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n476), .A2(G270), .A3(new_n289), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n586), .A2(new_n587), .A3(new_n475), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n586), .B2(new_n475), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n580), .A2(G169), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G179), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n580), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n566), .A2(new_n568), .A3(new_n565), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n572), .A2(new_n573), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n563), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n576), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n599), .A2(new_n600), .A3(new_n578), .ZN(new_n601));
  OAI211_X1 g0401(.A(G190), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n586), .A2(new_n475), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT85), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n586), .A2(new_n587), .A3(new_n475), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n604), .A2(new_n605), .B1(new_n582), .B2(new_n584), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n601), .B(new_n602), .C1(new_n515), .C2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n580), .A2(KEYINPUT21), .A3(G169), .A4(new_n590), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n593), .A2(new_n596), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n357), .A2(new_n223), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n511), .B2(new_n223), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n323), .A2(G97), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n223), .A2(G107), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g0415(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT78), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(KEYINPUT6), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT6), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(KEYINPUT78), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n613), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n622), .A3(G20), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT79), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n258), .A2(G77), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n323), .B1(new_n414), .B2(new_n415), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n612), .B1(new_n629), .B2(new_n342), .ZN(new_n630));
  INV_X1    g0430(.A(new_n567), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n283), .A2(new_n285), .A3(G244), .A4(new_n280), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT4), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n283), .A2(new_n285), .A3(G250), .A4(G1698), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT80), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT80), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n279), .A2(new_n638), .A3(G250), .A4(G1698), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n634), .A2(new_n635), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n290), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n476), .A2(G257), .A3(new_n289), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n475), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(G169), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  AOI211_X1 g0445(.A(G179), .B(new_n643), .C1(new_n640), .C2(new_n290), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n630), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n623), .A2(new_n625), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT79), .ZN(new_n650));
  INV_X1    g0450(.A(new_n628), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n611), .B1(new_n653), .B2(new_n252), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n641), .A2(new_n644), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G200), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n643), .B1(new_n640), .B2(new_n290), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G190), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n560), .A2(new_n609), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n461), .A2(new_n661), .ZN(G372));
  NAND2_X1  g0462(.A1(new_n479), .A2(new_n481), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n501), .B2(new_n512), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n593), .A2(new_n664), .A3(new_n596), .A4(new_n608), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT90), .B1(new_n532), .B2(new_n515), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT90), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(G200), .C1(new_n535), .C2(new_n523), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n558), .A2(new_n666), .A3(new_n553), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n532), .A2(new_n533), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n540), .A2(new_n551), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n514), .B2(new_n517), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n665), .A2(new_n673), .A3(new_n648), .A4(new_n659), .ZN(new_n674));
  INV_X1    g0474(.A(new_n671), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n657), .A2(new_n533), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(G169), .B2(new_n657), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n672), .A2(new_n677), .A3(new_n654), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n677), .A2(new_n654), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n559), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n674), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n461), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n388), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n312), .A2(new_n273), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n345), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n302), .A3(new_n458), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n459), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n686), .B1(new_n690), .B2(new_n382), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n593), .A2(new_n596), .A3(new_n608), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n356), .A2(G20), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n275), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n601), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n609), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n499), .B1(new_n498), .B2(new_n492), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n252), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n511), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n506), .A2(new_n508), .B1(new_n710), .B2(G107), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n706), .A2(new_n482), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n709), .A2(new_n711), .A3(new_n517), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n514), .B2(new_n701), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n513), .B2(new_n701), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n705), .A2(G330), .A3(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n664), .A2(new_n700), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n693), .A2(new_n701), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n714), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n209), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n542), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n233), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n724), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(G330), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n513), .A2(new_n518), .A3(new_n559), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n596), .A2(new_n593), .A3(new_n608), .A4(new_n607), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n648), .A2(new_n659), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n701), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n655), .A2(KEYINPUT92), .A3(new_n478), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n539), .A2(new_n533), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n606), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT92), .ZN(new_n739));
  INV_X1    g0539(.A(new_n478), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n657), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n736), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n604), .A2(new_n605), .ZN(new_n744));
  INV_X1    g0544(.A(new_n477), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n289), .B1(new_n464), .B2(new_n465), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n744), .A2(G179), .A3(new_n585), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n657), .A2(new_n532), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n641), .A2(new_n644), .A3(new_n532), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(new_n595), .A3(KEYINPUT30), .A4(new_n747), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n742), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n700), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT93), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT93), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n753), .A2(new_n758), .A3(KEYINPUT31), .A4(new_n700), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n730), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n684), .A2(new_n701), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n513), .A2(new_n596), .A3(new_n608), .A4(new_n593), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT94), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n648), .A2(new_n659), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(new_n648), .B2(new_n659), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n673), .B(new_n766), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(KEYINPUT26), .B1(new_n648), .B2(new_n672), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n681), .A2(new_n559), .A3(new_n679), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n770), .A2(new_n671), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(KEYINPUT29), .A3(new_n701), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n762), .B1(new_n765), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n729), .B1(new_n775), .B2(G1), .ZN(G364));
  NAND2_X1  g0576(.A1(new_n694), .A2(G45), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n724), .A2(G1), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n705), .B2(G330), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G330), .B2(new_n705), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n228), .B1(G20), .B2(new_n307), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n229), .A2(new_n533), .A3(new_n347), .A4(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n318), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT98), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n515), .B2(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n533), .A2(KEYINPUT98), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n229), .A2(G190), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G179), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G329), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n792), .A2(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n229), .B1(new_n794), .B2(G190), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(G294), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n229), .A2(new_n347), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n789), .A2(new_n801), .A3(new_n790), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n800), .B1(new_n583), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n533), .A2(new_n515), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n804), .A2(new_n791), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n787), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n347), .A2(new_n515), .A3(G20), .A4(G179), .ZN(new_n809));
  INV_X1    g0609(.A(G326), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n804), .A2(new_n801), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT99), .Z(new_n812));
  OAI221_X1 g0612(.A(new_n807), .B1(new_n808), .B2(new_n809), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n792), .A2(new_n323), .ZN(new_n814));
  INV_X1    g0614(.A(new_n802), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G87), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n795), .A2(new_n402), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n279), .B1(new_n785), .B2(new_n202), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n811), .A2(new_n232), .B1(new_n798), .B2(new_n223), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(new_n817), .C2(new_n819), .ZN(new_n824));
  INV_X1    g0624(.A(new_n805), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n203), .B2(new_n825), .C1(new_n263), .C2(new_n809), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n783), .B1(new_n813), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(G13), .A2(G33), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(G20), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n782), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT96), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n279), .A2(G355), .A3(new_n209), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n246), .A2(G45), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n722), .A2(new_n279), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n727), .B2(G45), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n833), .B1(G116), .B2(new_n209), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n827), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n778), .B(KEYINPUT95), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n830), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n838), .B(new_n840), .C1(new_n704), .C2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n781), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  OAI22_X1  g0644(.A1(new_n808), .A2(new_n795), .B1(new_n798), .B2(new_n223), .ZN(new_n845));
  INV_X1    g0645(.A(new_n811), .ZN(new_n846));
  INV_X1    g0646(.A(new_n809), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n846), .A2(G303), .B1(new_n494), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n793), .B2(new_n825), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT100), .Z(new_n850));
  INV_X1    g0650(.A(new_n792), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n845), .B(new_n850), .C1(G87), .C2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n318), .B1(new_n802), .B2(new_n323), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT101), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n852), .B(new_n854), .C1(new_n855), .C2(new_n785), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT102), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G150), .A2(new_n805), .B1(new_n784), .B2(G143), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n811), .C1(new_n402), .C2(new_n809), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n851), .A2(G68), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n815), .A2(G50), .B1(G58), .B2(new_n799), .ZN(new_n863));
  INV_X1    g0663(.A(new_n795), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n318), .B1(new_n864), .B2(G132), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n783), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n782), .A2(new_n828), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n839), .B(new_n867), .C1(new_n263), .C2(new_n868), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n329), .A2(new_n343), .A3(new_n344), .A4(new_n701), .ZN(new_n870));
  INV_X1    g0670(.A(new_n345), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n348), .A2(new_n349), .B1(new_n343), .B2(new_n700), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n829), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n684), .A2(new_n351), .A3(new_n701), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n763), .B2(new_n873), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(new_n762), .Z(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n778), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(G384));
  NAND2_X1  g0681(.A1(new_n273), .A2(new_n700), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n687), .A2(new_n302), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n312), .A2(new_n273), .A3(new_n700), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n876), .A2(new_n870), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n398), .B2(new_n405), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n408), .B2(new_n409), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n394), .B1(new_n888), .B2(new_n257), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n452), .B1(new_n430), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n698), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n698), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n438), .A2(new_n394), .B1(new_n429), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n452), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n891), .B1(new_n440), .B2(new_n456), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n885), .B(new_n886), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n459), .A2(new_n893), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT103), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n421), .A2(new_n698), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n440), .B2(new_n456), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n894), .A2(new_n452), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n896), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n687), .A2(new_n700), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n888), .A2(new_n257), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n893), .B1(new_n919), .B2(new_n394), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n458), .B2(new_n459), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n894), .A2(new_n895), .A3(new_n452), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n429), .B1(new_n919), .B2(new_n394), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n923), .A3(new_n452), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n912), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n917), .A2(new_n918), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT103), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n901), .A2(new_n929), .A3(new_n903), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n905), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n774), .A2(new_n461), .A3(new_n765), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n691), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n931), .B(new_n933), .Z(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n756), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT31), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n661), .B2(new_n701), .ZN(new_n938));
  INV_X1    g0738(.A(new_n754), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n734), .B2(KEYINPUT31), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n756), .B(KEYINPUT104), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT105), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n941), .B1(KEYINPUT105), .B2(KEYINPUT40), .C1(new_n942), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n926), .A2(new_n914), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  INV_X1    g0750(.A(new_n944), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n915), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n461), .B(new_n940), .C1(new_n949), .C2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n944), .A2(new_n945), .B1(new_n926), .B2(new_n914), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n907), .B2(new_n910), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n940), .B(new_n941), .C1(new_n899), .C2(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n954), .A2(new_n947), .B1(new_n956), .B2(KEYINPUT40), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n730), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n461), .A2(new_n940), .A3(G330), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n953), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n934), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n275), .B2(new_n694), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n617), .A2(new_n622), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT35), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n229), .B(new_n228), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n966), .B(G116), .C1(new_n965), .C2(new_n964), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT36), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n233), .A2(G77), .A3(new_n399), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(G50), .B2(new_n203), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(G1), .A3(new_n356), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n963), .A2(new_n968), .A3(new_n971), .ZN(G367));
  OR2_X1    g0772(.A1(new_n768), .A2(new_n769), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(new_n714), .A3(new_n719), .A4(new_n766), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT42), .Z(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(new_n654), .B2(new_n701), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n648), .B1(new_n976), .B2(new_n513), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n701), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n701), .A2(new_n558), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n675), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n672), .B2(new_n980), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n979), .A2(KEYINPUT43), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT106), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n982), .B(KEYINPUT43), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT107), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n988), .A3(KEYINPUT108), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT108), .B1(new_n985), .B2(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n681), .A2(new_n700), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n976), .A2(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n990), .A2(new_n991), .B1(new_n717), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n991), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n717), .A2(new_n993), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n996), .A3(new_n989), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n723), .B(KEYINPUT41), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n720), .A2(new_n718), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT44), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n993), .A2(new_n1000), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n717), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n705), .A2(G330), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT109), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n720), .B1(new_n716), .B2(new_n719), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n775), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n999), .B1(new_n1011), .B2(new_n775), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n777), .A2(G1), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n994), .B(new_n997), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n812), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(G143), .B1(G68), .B2(new_n799), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n353), .B2(new_n785), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT111), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n805), .A2(G159), .B1(new_n847), .B2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n318), .B(new_n1020), .C1(G58), .C2(new_n815), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n851), .A2(G77), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n795), .A2(new_n859), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT46), .B1(new_n815), .B2(new_n494), .ZN(new_n1025));
  INV_X1    g0825(.A(G317), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n318), .B1(new_n795), .B2(new_n1026), .C1(new_n792), .C2(new_n223), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT110), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1025), .B(new_n1029), .C1(G294), .C2(new_n805), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n784), .A2(G303), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n815), .A2(KEYINPUT46), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G116), .A2(new_n1032), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1015), .A2(G311), .B1(G283), .B2(new_n847), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n798), .A2(new_n323), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1023), .A2(new_n1024), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT47), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n782), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n982), .A2(new_n841), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n835), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n831), .B1(new_n209), .B2(new_n339), .C1(new_n242), .C2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1039), .A2(new_n840), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1014), .A2(new_n1043), .ZN(G387));
  OAI21_X1  g0844(.A(new_n318), .B1(new_n795), .B2(new_n810), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n815), .A2(G294), .B1(G283), .B2(new_n799), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n805), .B1(new_n784), .B2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n583), .B2(new_n809), .C1(new_n812), .C2(new_n786), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT115), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT49), .Z(new_n1054));
  AOI211_X1 g0854(.A(new_n1045), .B(new_n1054), .C1(new_n494), .C2(new_n851), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n802), .A2(new_n263), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n223), .B2(new_n792), .C1(new_n353), .C2(new_n795), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n550), .A2(new_n798), .B1(new_n333), .B2(new_n825), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n785), .A2(new_n232), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n279), .B1(new_n203), .B2(new_n809), .C1(new_n811), .C2(new_n402), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n782), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n716), .A2(new_n841), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n725), .B(new_n473), .C1(new_n203), .C2(new_n263), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT113), .Z(new_n1066));
  OR3_X1    g0866(.A1(new_n333), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT50), .B1(new_n333), .B2(G50), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n239), .A2(G45), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n835), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n279), .A2(new_n209), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(G107), .B2(new_n209), .C1(new_n725), .C2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT114), .Z(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n832), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1063), .A2(new_n840), .A3(new_n1064), .A4(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1010), .A2(new_n775), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1010), .A2(new_n775), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n723), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1081), .ZN(G393));
  NAND2_X1  g0882(.A1(new_n993), .A2(new_n830), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n279), .B1(new_n333), .B2(new_n809), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n825), .A2(new_n232), .B1(new_n798), .B2(new_n263), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G87), .C2(new_n851), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n785), .A2(new_n402), .B1(new_n811), .B2(new_n353), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n864), .A2(G143), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n815), .A2(G68), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n318), .B1(new_n795), .B2(new_n786), .C1(new_n493), .C2(new_n798), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n814), .B(new_n1092), .C1(G303), .C2(new_n805), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n785), .A2(new_n808), .B1(new_n811), .B2(new_n1026), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT52), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n793), .C2(new_n802), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n809), .A2(new_n855), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n782), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n831), .B1(new_n223), .B2(new_n209), .C1(new_n249), .C2(new_n1041), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1083), .A2(new_n840), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1006), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1013), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n724), .B1(new_n1102), .B2(new_n1080), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1011), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  INV_X1    g0907(.A(KEYINPUT117), .ZN(new_n1108));
  OAI211_X1 g0908(.A(G330), .B(new_n874), .C1(new_n942), .C2(new_n760), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n883), .A2(new_n884), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n940), .A2(G330), .A3(new_n941), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n886), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n755), .A2(new_n761), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1115), .A2(G330), .A3(new_n874), .A4(new_n885), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n874), .C1(new_n942), .C2(new_n943), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1110), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n773), .A2(new_n351), .A3(new_n701), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n870), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n932), .A2(new_n959), .A3(new_n691), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1108), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(KEYINPUT117), .B(new_n1122), .C1(new_n1114), .C2(new_n1120), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n918), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n886), .A2(new_n885), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n917), .A2(new_n927), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n915), .A2(new_n1127), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1110), .B1(new_n1119), .B2(new_n870), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1112), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n927), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT39), .B1(new_n913), .B2(new_n914), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1110), .B1(new_n876), .B2(new_n870), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1134), .A2(new_n1135), .B1(new_n918), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1131), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n915), .A3(new_n1127), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1116), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1126), .A2(new_n1133), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1133), .A2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n723), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n828), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  AND2_X1   g0947(.A1(new_n1147), .A2(new_n847), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n815), .A2(G150), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n318), .B(new_n1148), .C1(new_n1149), .C2(KEYINPUT53), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n795), .C1(new_n1152), .C2(new_n811), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n798), .A2(new_n402), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n825), .A2(new_n859), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n851), .A2(G50), .B1(new_n784), .B2(G132), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(KEYINPUT53), .B2(new_n1149), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n815), .A2(G87), .B1(new_n846), .B2(G283), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n862), .C1(new_n220), .C2(new_n785), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n809), .A2(new_n223), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n825), .A2(new_n323), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n318), .B1(new_n798), .B2(new_n263), .C1(new_n855), .C2(new_n795), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n782), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n840), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n333), .B2(new_n868), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1143), .A2(new_n1013), .B1(new_n1146), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1145), .A2(new_n1168), .ZN(G378));
  INV_X1    g0969(.A(KEYINPUT122), .ZN(new_n1170));
  AOI211_X1 g0970(.A(KEYINPUT103), .B(new_n902), .C1(new_n948), .C2(new_n1136), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n929), .B1(new_n901), .B2(new_n903), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1170), .B1(new_n1173), .B2(new_n928), .ZN(new_n1174));
  AND4_X1   g0974(.A1(new_n1170), .A2(new_n905), .A3(new_n928), .A4(new_n930), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT120), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n382), .A2(new_n388), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n361), .A2(new_n893), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1183), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n958), .A2(new_n1177), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT120), .B1(new_n957), .B2(new_n730), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1177), .B(G330), .C1(new_n949), .C2(new_n952), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1188), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1176), .A2(KEYINPUT121), .A3(new_n1190), .A4(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(KEYINPUT121), .A3(new_n1190), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n931), .B(KEYINPUT122), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1144), .A2(new_n1123), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT123), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT123), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1203), .A3(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1193), .A2(new_n1190), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(new_n931), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n931), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1198), .A4(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1202), .A2(new_n723), .A3(new_n1204), .A4(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1194), .A2(new_n1197), .A3(new_n1013), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1189), .A2(new_n828), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1056), .B1(G116), .B2(new_n846), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n318), .C1(new_n202), .C2(new_n792), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n471), .B1(new_n203), .B2(new_n798), .C1(new_n550), .C2(new_n809), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G107), .C2(new_n784), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n223), .B2(new_n825), .C1(new_n793), .C2(new_n795), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n815), .A2(new_n1147), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(KEYINPUT118), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(KEYINPUT118), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n805), .A2(G132), .B1(new_n847), .B2(G137), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1220), .B(new_n1223), .C1(G128), .C2(new_n784), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n1151), .B2(new_n811), .C1(new_n353), .C2(new_n798), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G41), .B1(new_n1225), .B2(KEYINPUT59), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G33), .B1(new_n864), .B2(G124), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n402), .C2(new_n792), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1217), .B1(G50), .B2(new_n1218), .C1(new_n1226), .C2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT119), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n782), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n868), .A2(new_n232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1211), .A2(new_n1232), .A3(new_n779), .A4(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1210), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1209), .A2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1121), .A2(new_n1013), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n550), .A2(new_n798), .B1(new_n855), .B2(new_n811), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1022), .B1(new_n223), .B2(new_n802), .C1(new_n793), .C2(new_n785), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n318), .B1(new_n809), .B2(new_n323), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n583), .B2(new_n795), .C1(new_n493), .C2(new_n825), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G58), .A2(new_n851), .B1(new_n846), .B2(G132), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n1152), .B2(new_n795), .C1(new_n402), .C2(new_n802), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G137), .B2(new_n784), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n805), .A2(new_n1147), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n799), .A2(G50), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n318), .B1(new_n847), .B2(G150), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n783), .B1(new_n1242), .B2(new_n1249), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n839), .B(new_n1250), .C1(new_n203), .C2(new_n868), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n885), .B2(new_n829), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1237), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1114), .A2(new_n1122), .A3(new_n1120), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1126), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1256), .B2(new_n999), .ZN(G381));
  XNOR2_X1  g1057(.A(G378), .B(KEYINPUT124), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G375), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G384), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(G393), .A2(G381), .A3(G396), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1014), .A2(new_n1043), .A3(new_n1106), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1264), .ZN(G407));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1260), .B2(new_n699), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(G407), .ZN(G409));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1255), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1256), .B2(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n723), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1254), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(G384), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1266), .A2(G343), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(G2897), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT126), .Z(new_n1277));
  XNOR2_X1  g1077(.A(new_n1274), .B(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1209), .A2(G378), .A3(new_n1235), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1206), .A2(new_n1013), .A3(new_n1207), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1280), .B(new_n1234), .C1(new_n1199), .C2(new_n999), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1258), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1275), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(new_n843), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1106), .B1(new_n1014), .B2(new_n1043), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1264), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(G390), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1287), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1263), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1273), .B(new_n1261), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n1275), .B(new_n1294), .C1(new_n1279), .C2(new_n1282), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1295), .B2(KEYINPUT63), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1283), .A2(new_n1298), .A3(new_n1284), .A4(new_n1274), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1286), .B(new_n1296), .C1(new_n1299), .C2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT62), .B1(new_n1300), .B2(KEYINPUT127), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1294), .B(new_n1277), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1275), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT125), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1306), .B2(new_n1274), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1303), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1264), .A2(new_n1288), .A3(new_n1287), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1291), .B1(new_n1290), .B2(new_n1263), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1302), .B1(new_n1310), .B2(new_n1313), .ZN(G405));
  INV_X1    g1114(.A(new_n1279), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1259), .B1(new_n1235), .B2(new_n1209), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1293), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1294), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1317), .A2(new_n1274), .A3(new_n1319), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


