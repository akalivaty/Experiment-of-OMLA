//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n217), .B1(KEYINPUT67), .B2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n209), .B(new_n220), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G33), .A3(G41), .ZN(new_n254));
  INV_X1    g0054(.A(new_n221), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n248), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n250), .B1(new_n258), .B2(G238), .ZN(new_n259));
  INV_X1    g0059(.A(new_n251), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT70), .B1(new_n225), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT70), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(new_n251), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G226), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G97), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT76), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n267), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n267), .B2(new_n273), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n259), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n279), .B(new_n259), .C1(new_n275), .C2(new_n276), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n278), .A2(KEYINPUT77), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT77), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n277), .A2(new_n282), .A3(KEYINPUT13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(G179), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  AOI211_X1 g0086(.A(KEYINPUT14), .B(new_n286), .C1(new_n278), .C2(new_n280), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n278), .A2(new_n280), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT14), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(G77), .B1(G20), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n202), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT71), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n225), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n226), .A2(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G13), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n295), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT12), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n305), .A2(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G68), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n292), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(G190), .B1(new_n281), .B2(new_n284), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n289), .B2(G200), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT78), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT78), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n314), .A2(G77), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n311), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n329), .A2(new_n298), .B1(new_n226), .B2(new_n327), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT15), .B(G87), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n226), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n305), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n326), .A2(new_n328), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n250), .B1(new_n258), .B2(G244), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n293), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G232), .ZN(new_n344));
  INV_X1    g0144(.A(G107), .ZN(new_n345));
  INV_X1    g0145(.A(G238), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n268), .A2(G1698), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n344), .B1(new_n345), .B2(new_n268), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n338), .B1(new_n348), .B2(new_n267), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n336), .B1(new_n350), .B2(new_n286), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(new_n349), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT75), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n358), .A2(KEYINPUT75), .B1(G190), .B2(new_n349), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n354), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n302), .A2(new_n303), .B1(new_n223), .B2(new_n224), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n329), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n294), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n314), .A2(G50), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n311), .A2(new_n202), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n343), .A2(G222), .ZN(new_n372));
  INV_X1    g0172(.A(G223), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n372), .B1(new_n327), .B2(new_n268), .C1(new_n373), .C2(new_n347), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n267), .ZN(new_n375));
  INV_X1    g0175(.A(new_n250), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n257), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT69), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n382), .B2(new_n286), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G179), .B2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT73), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(KEYINPUT73), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n361), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n371), .A2(KEYINPUT9), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT9), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n367), .B2(new_n370), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n388), .B(new_n390), .C1(new_n391), .C2(new_n382), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n382), .A2(G200), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n388), .A2(new_n390), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT10), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n382), .A2(new_n391), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n393), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n268), .A2(new_n270), .ZN(new_n401));
  INV_X1    g0201(.A(G87), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n401), .A2(new_n373), .B1(new_n293), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n347), .A2(new_n377), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n267), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n250), .B1(new_n258), .B2(G232), .ZN(new_n406));
  AOI21_X1  g0206(.A(G169), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n409), .B2(new_n352), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n268), .A2(new_n411), .A3(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n342), .B2(new_n226), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n297), .A2(G159), .ZN(new_n415));
  INV_X1    g0215(.A(G58), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n295), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n417), .B2(new_n201), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n411), .B1(new_n268), .B2(G20), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n295), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n415), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n305), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n364), .A2(new_n310), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n314), .B2(new_n364), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT18), .B1(new_n410), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n410), .A2(KEYINPUT18), .A3(new_n429), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n408), .A2(G200), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n405), .A2(G190), .A3(new_n406), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n426), .A3(new_n428), .A4(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n400), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n387), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n323), .A2(new_n325), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n298), .A2(new_n327), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n345), .A2(G97), .ZN(new_n442));
  INV_X1    g0242(.A(G97), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G107), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n445), .B2(new_n442), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n441), .B1(new_n447), .B2(G20), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n345), .B1(new_n421), .B2(new_n422), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT79), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI211_X1 g0251(.A(KEYINPUT79), .B(new_n345), .C1(new_n421), .C2(new_n422), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n305), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n310), .A2(G97), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n309), .A2(G13), .B1(new_n247), .B2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n304), .A3(new_n225), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n362), .A2(KEYINPUT80), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n454), .B1(new_n460), .B2(G97), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(new_n270), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n270), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n267), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n471), .A2(new_n473), .A3(new_n247), .A4(G45), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n256), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n473), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n247), .A2(G45), .A3(G274), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n478), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(KEYINPUT82), .A3(new_n471), .A4(new_n473), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n475), .A2(G257), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n469), .A2(G190), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n453), .A2(new_n461), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n267), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT81), .B1(new_n468), .B2(new_n267), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G200), .ZN(new_n488));
  AOI21_X1  g0288(.A(G169), .B1(new_n469), .B2(new_n482), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n453), .B2(new_n461), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n352), .B(new_n482), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n484), .A2(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n331), .B1(new_n458), .B2(new_n459), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n226), .B1(new_n272), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n402), .A2(new_n443), .A3(new_n345), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n339), .A2(new_n341), .A3(new_n226), .A4(G68), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n332), .B2(new_n443), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n305), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n311), .A2(new_n331), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT85), .B1(new_n493), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n331), .ZN(new_n505));
  AND4_X1   g0305(.A1(KEYINPUT80), .A2(new_n455), .A3(new_n304), .A4(new_n225), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT80), .B1(new_n362), .B2(new_n455), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n500), .A2(new_n305), .B1(new_n311), .B2(new_n331), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n339), .A2(new_n341), .A3(G238), .A4(new_n270), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT84), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT84), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G116), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n518), .A3(G33), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n265), .B1(new_n264), .B2(new_n251), .ZN(new_n521));
  AND4_X1   g0321(.A1(new_n265), .A2(new_n223), .A3(new_n224), .A4(new_n251), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  INV_X1    g0324(.A(G45), .ZN(new_n525));
  OAI21_X1  g0325(.A(G250), .B1(new_n525), .B2(G1), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n256), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n528), .B2(new_n478), .ZN(new_n529));
  AOI211_X1 g0329(.A(KEYINPUT83), .B(new_n480), .C1(new_n256), .C2(new_n527), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n523), .B(new_n352), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n221), .B1(KEYINPUT68), .B2(new_n251), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n526), .B1(new_n533), .B2(new_n254), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT83), .B1(new_n534), .B2(new_n480), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n528), .A2(new_n524), .A3(new_n478), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(G169), .B1(new_n537), .B2(new_n523), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(G87), .B1(new_n506), .B2(new_n507), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n510), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n357), .B1(new_n537), .B2(new_n523), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n535), .A2(new_n536), .B1(new_n267), .B2(new_n520), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n512), .A2(new_n539), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n339), .A2(new_n341), .A3(new_n226), .A4(G87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n268), .A2(new_n549), .A3(new_n226), .A4(G87), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n226), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n345), .A2(KEYINPUT23), .A3(G20), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n294), .A2(new_n516), .A3(new_n518), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT24), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n548), .B2(new_n550), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT86), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n305), .ZN(new_n567));
  OAI21_X1  g0367(.A(G107), .B1(new_n506), .B2(new_n507), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n311), .A2(new_n345), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(KEYINPUT87), .A3(KEYINPUT25), .ZN(new_n570));
  XNOR2_X1  g0370(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n339), .A2(new_n341), .A3(G250), .A4(new_n270), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(G1698), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(new_n576), .C1(new_n293), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n267), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n479), .A2(new_n481), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n475), .A2(G264), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n357), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n267), .A2(new_n578), .B1(new_n475), .B2(G264), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n391), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AND4_X1   g0386(.A1(KEYINPUT89), .A2(new_n567), .A3(new_n574), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n573), .B1(new_n566), .B2(new_n305), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT89), .B1(new_n588), .B2(new_n586), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n492), .B(new_n546), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n567), .A2(new_n574), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(new_n286), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n584), .A2(new_n352), .A3(new_n580), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(KEYINPUT88), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n593), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n516), .A2(new_n518), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G20), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n467), .B(new_n226), .C1(G33), .C2(new_n443), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n305), .A2(KEYINPUT20), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g0405(.A(KEYINPUT84), .B(G116), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(new_n226), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n607), .B2(new_n362), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n311), .A2(new_n601), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n362), .A2(G116), .A3(new_n455), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n475), .A2(G270), .B1(new_n479), .B2(new_n481), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(new_n270), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n339), .A2(new_n341), .A3(G264), .A4(G1698), .ZN(new_n615));
  INV_X1    g0415(.A(G303), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n268), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n267), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n286), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT21), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n612), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n613), .A2(new_n618), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n613), .A2(new_n618), .A3(G190), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n612), .A2(new_n619), .A3(KEYINPUT21), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n256), .A2(new_n474), .A3(G270), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n580), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n267), .B2(new_n617), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n612), .A2(new_n630), .A3(G179), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n621), .A2(new_n626), .A3(new_n627), .A4(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n440), .A2(new_n590), .A3(new_n600), .A4(new_n632), .ZN(G372));
  AND3_X1   g0433(.A1(new_n323), .A2(new_n325), .A3(new_n439), .ZN(new_n634));
  INV_X1    g0434(.A(new_n489), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n345), .A2(KEYINPUT6), .A3(G97), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n244), .B2(new_n445), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n637), .A2(new_n226), .B1(new_n327), .B2(new_n298), .ZN(new_n638));
  OAI21_X1  g0438(.A(G107), .B1(new_n412), .B2(new_n413), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(KEYINPUT79), .ZN(new_n640));
  INV_X1    g0440(.A(new_n452), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n362), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n460), .A2(G97), .ZN(new_n643));
  INV_X1    g0443(.A(new_n454), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n635), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n491), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT81), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n469), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n267), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n357), .B1(new_n651), .B2(new_n482), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n453), .A2(new_n461), .A3(new_n483), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n646), .A2(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n503), .B1(G87), .B2(new_n460), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n545), .B(new_n655), .C1(new_n357), .C2(new_n544), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n493), .A2(new_n503), .A3(KEYINPUT85), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n531), .B1(new_n544), .B2(G169), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n551), .A2(new_n563), .A3(new_n558), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n563), .B1(new_n551), .B2(new_n558), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n560), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n362), .B1(new_n666), .B2(new_n564), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n663), .B(new_n594), .C1(new_n667), .C2(new_n573), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT90), .B1(new_n588), .B2(new_n597), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n627), .A2(new_n631), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n620), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n567), .A2(new_n586), .A3(new_n574), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT89), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n588), .A2(KEYINPUT89), .A3(new_n586), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n662), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n512), .A2(new_n539), .A3(KEYINPUT91), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT91), .B1(new_n512), .B2(new_n539), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n490), .A2(new_n491), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n661), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n453), .A2(new_n461), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n685), .A2(new_n491), .A3(new_n635), .ZN(new_n686));
  XOR2_X1   g0486(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n687));
  NAND3_X1  g0487(.A1(new_n546), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n681), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n634), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n386), .A2(new_n385), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n354), .B1(new_n292), .B2(new_n317), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n321), .A2(new_n437), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n433), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n695), .B2(new_n400), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(G369));
  AND2_X1   g0497(.A1(new_n226), .A2(G13), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n247), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n677), .B(new_n599), .C1(new_n588), .C2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n591), .A2(new_n594), .A3(new_n704), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n621), .A2(new_n627), .A3(new_n631), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n622), .A2(new_n705), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n632), .B2(new_n711), .ZN(new_n713));
  XNOR2_X1  g0513(.A(KEYINPUT93), .B(G330), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n599), .A2(new_n677), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n710), .A2(new_n705), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n668), .A2(new_n669), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n705), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0524(.A(new_n207), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n496), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n229), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n710), .B1(new_n595), .B2(new_n598), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n590), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n679), .A2(new_n680), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n546), .A2(new_n686), .A3(new_n682), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n687), .B1(new_n661), .B2(new_n683), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n705), .C1(new_n733), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n704), .B1(new_n678), .B2(new_n689), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(KEYINPUT29), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n714), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n630), .A2(G179), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n742), .A2(new_n487), .A3(new_n582), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n544), .A2(G179), .A3(new_n618), .A4(new_n613), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n584), .A2(new_n482), .A3(new_n469), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT95), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n623), .A2(new_n743), .A3(new_n352), .ZN(new_n752));
  INV_X1    g0552(.A(new_n747), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(KEYINPUT30), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n744), .A2(KEYINPUT95), .A3(new_n748), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT31), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n705), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n744), .A2(new_n754), .A3(new_n748), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n704), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n756), .A2(new_n758), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n632), .B1(new_n595), .B2(new_n598), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(new_n662), .A3(new_n677), .A4(new_n705), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n741), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n740), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n731), .B1(new_n767), .B2(G1), .ZN(G364));
  AOI21_X1  g0568(.A(new_n247), .B1(new_n698), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n726), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n713), .B2(new_n714), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n714), .B2(new_n713), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n725), .A2(new_n342), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G355), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G116), .B2(new_n207), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n242), .A2(new_n525), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n725), .A2(new_n268), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n525), .B2(new_n230), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n783), .A2(KEYINPUT96), .A3(G20), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT96), .B1(new_n783), .B2(G20), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n225), .B1(G20), .B2(new_n286), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n771), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n226), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n357), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n352), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n791), .A2(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n352), .A2(new_n357), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n792), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G317), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(KEYINPUT33), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n226), .A2(new_n391), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n795), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n799), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n798), .B(new_n809), .C1(G326), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G179), .A2(G200), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  INV_X1    g0614(.A(new_n792), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G329), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n807), .A2(new_n793), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n342), .B1(new_n818), .B2(new_n616), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  OAI21_X1  g0620(.A(G20), .B1(new_n814), .B2(new_n391), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G294), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n812), .A2(new_n817), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n816), .A2(G159), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT32), .Z(new_n825));
  INV_X1    g0625(.A(new_n796), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n811), .A2(G50), .B1(new_n826), .B2(G77), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n295), .B2(new_n800), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n268), .B1(new_n794), .B2(new_n345), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n416), .A2(new_n808), .B1(new_n818), .B2(new_n402), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n821), .A2(G97), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n825), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n790), .B1(new_n834), .B2(new_n787), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n786), .B(KEYINPUT99), .Z(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n713), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n773), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  INV_X1    g0639(.A(new_n771), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n787), .A2(new_n782), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n327), .ZN(new_n842));
  INV_X1    g0642(.A(new_n787), .ZN(new_n843));
  INV_X1    g0643(.A(new_n808), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G283), .A2(new_n801), .B1(new_n844), .B2(G294), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n345), .B2(new_n818), .ZN(new_n846));
  INV_X1    g0646(.A(new_n794), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G87), .A2(new_n847), .B1(new_n826), .B2(new_n606), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n342), .C1(new_n616), .C2(new_n810), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n846), .B(new_n849), .C1(G311), .C2(new_n816), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n794), .A2(new_n295), .ZN(new_n851));
  INV_X1    g0651(.A(new_n818), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n342), .B(new_n851), .C1(G50), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  INV_X1    g0654(.A(new_n816), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n857), .A2(new_n808), .B1(new_n800), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  INV_X1    g0660(.A(G159), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n810), .A2(new_n860), .B1(new_n796), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n856), .B1(KEYINPUT34), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G58), .B2(new_n821), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n832), .A2(new_n850), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n354), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n704), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n359), .A2(new_n360), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n336), .B2(new_n705), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n871), .B2(new_n868), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n842), .B1(new_n843), .B2(new_n867), .C1(new_n872), .C2(new_n783), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT100), .ZN(new_n874));
  AND4_X1   g0674(.A1(new_n874), .A2(new_n690), .A3(new_n361), .A4(new_n705), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n739), .B2(new_n361), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n875), .A2(new_n876), .B1(new_n739), .B2(new_n872), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n771), .B1(new_n877), .B2(new_n765), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n765), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(G384));
  OAI211_X1 g0681(.A(G116), .B(new_n227), .C1(new_n447), .C2(KEYINPUT35), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(KEYINPUT35), .B2(new_n447), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT36), .ZN(new_n884));
  OR3_X1    g0684(.A1(new_n229), .A2(new_n327), .A3(new_n417), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n202), .A2(G68), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n247), .B(G13), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n317), .A2(new_n704), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n278), .A2(KEYINPUT77), .A3(new_n280), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n352), .B1(new_n890), .B2(new_n283), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT14), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n289), .B2(G169), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n891), .A2(new_n893), .A3(new_n287), .ZN(new_n894));
  INV_X1    g0694(.A(new_n317), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n321), .B(new_n889), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n292), .A2(new_n317), .A3(new_n704), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n757), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n760), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n759), .A2(new_n899), .A3(new_n757), .A4(new_n704), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n763), .A2(new_n903), .A3(KEYINPUT103), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT103), .B1(new_n763), .B2(new_n903), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n898), .B(new_n872), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n410), .A2(new_n429), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n702), .B1(new_n426), .B2(new_n428), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n910), .A3(new_n436), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n433), .B2(new_n437), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n432), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n430), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n909), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n909), .B2(KEYINPUT101), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n911), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n911), .A2(new_n922), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT40), .B1(new_n906), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n763), .A2(new_n903), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n763), .A2(new_n903), .A3(KEYINPUT103), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n924), .A2(new_n923), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n907), .B1(new_n933), .B2(new_n914), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT40), .B1(new_n934), .B2(new_n925), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n932), .A2(new_n935), .A3(new_n872), .A4(new_n898), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n634), .A2(new_n932), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n714), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n696), .B1(new_n440), .B2(new_n740), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n917), .A2(new_n702), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n915), .A2(new_n925), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n934), .B2(new_n925), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n318), .A2(new_n704), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n943), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n662), .A2(new_n672), .A3(new_n677), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n546), .A2(new_n686), .A3(new_n687), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT26), .B1(new_n546), .B2(new_n686), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n734), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n361), .B(new_n705), .C1(new_n952), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT100), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n739), .A2(new_n874), .A3(new_n361), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n869), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n898), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n934), .A2(new_n925), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n951), .A2(new_n963), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n942), .A2(new_n964), .B1(new_n247), .B2(new_n698), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n942), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n888), .B1(new_n965), .B2(new_n966), .ZN(G367));
  INV_X1    g0767(.A(KEYINPUT106), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n681), .A2(new_n541), .A3(new_n704), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT104), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(KEYINPUT104), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n546), .B1(new_n655), .B2(new_n705), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT43), .B1(new_n973), .B2(KEYINPUT105), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(KEYINPUT105), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n600), .B1(new_n652), .B2(new_n653), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n704), .B1(new_n976), .B2(new_n683), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT42), .ZN(new_n978));
  INV_X1    g0778(.A(new_n720), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n685), .A2(new_n704), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n492), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n686), .A2(new_n704), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n978), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n983), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n977), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n975), .B2(new_n987), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n968), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n975), .A2(new_n987), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n993), .A2(KEYINPUT106), .A3(new_n988), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n717), .A2(new_n984), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n726), .B(KEYINPUT41), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n709), .A2(new_n719), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n979), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n716), .B1(new_n1001), .B2(new_n715), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n767), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT107), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n722), .A2(new_n983), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(KEYINPUT44), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n722), .A2(new_n983), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT45), .B1(new_n722), .B2(new_n983), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1007), .A2(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n716), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n717), .B1(new_n1011), .B2(new_n1012), .C1(new_n1008), .C2(new_n1007), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT107), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1003), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1005), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n999), .B1(new_n1018), .B2(new_n767), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n997), .B1(new_n770), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT108), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n997), .B(KEYINPUT108), .C1(new_n770), .C2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n973), .A2(new_n836), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n788), .B1(new_n207), .B2(new_n331), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n238), .A2(new_n779), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n771), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT109), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G303), .A2(new_n844), .B1(new_n826), .B2(G283), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1030), .B(new_n342), .C1(new_n797), .C2(new_n810), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n852), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n443), .B2(new_n794), .C1(new_n577), .C2(new_n800), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n855), .A2(new_n802), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT46), .B1(new_n852), .B2(new_n606), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n821), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n345), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT110), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n810), .A2(new_n857), .B1(new_n796), .B2(new_n202), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n416), .A2(new_n818), .B1(new_n808), .B2(new_n858), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G159), .C2(new_n801), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n816), .A2(G137), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n268), .B1(new_n794), .B2(new_n327), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n821), .A2(G68), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT47), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n843), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1039), .A2(KEYINPUT47), .A3(new_n1047), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1029), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1025), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1024), .A2(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n1002), .A2(new_n770), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n779), .B1(new_n235), .B2(G45), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n728), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n774), .ZN(new_n1057));
  AOI21_X1  g0857(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n329), .A2(G50), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n728), .B(new_n1058), .C1(new_n1059), .C2(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT50), .B2(new_n1059), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1057), .A2(new_n1061), .B1(G107), .B2(new_n207), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n840), .B1(new_n1062), .B2(new_n788), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT112), .B(G150), .Z(new_n1064));
  AOI22_X1  g0864(.A1(new_n364), .A2(new_n801), .B1(new_n816), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n821), .A2(new_n505), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n810), .A2(new_n861), .B1(new_n808), .B2(new_n202), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n818), .A2(new_n327), .B1(new_n796), .B2(new_n295), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n268), .B1(new_n794), .B2(new_n443), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1065), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n811), .A2(G322), .B1(new_n826), .B2(G303), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n797), .B2(new_n800), .C1(new_n802), .C2(new_n808), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT113), .Z(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT48), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT48), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n821), .A2(G283), .B1(G294), .B2(new_n852), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT49), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n816), .A2(G326), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n342), .C1(new_n601), .C2(new_n794), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1071), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1063), .B1(new_n708), .B2(new_n836), .C1(new_n1084), .C2(new_n843), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1004), .A2(new_n727), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1086), .A2(KEYINPUT114), .B1(new_n767), .B2(new_n1002), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1054), .B(new_n1085), .C1(new_n1087), .C2(new_n1088), .ZN(G393));
  NAND2_X1  g0889(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1018), .B(new_n726), .C1(new_n1091), .C2(new_n1004), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n770), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n788), .B1(new_n443), .B2(new_n207), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n245), .A2(new_n779), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n771), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n810), .A2(new_n802), .B1(new_n808), .B2(new_n797), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT52), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n806), .C2(new_n855), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n800), .A2(new_n616), .B1(new_n796), .B2(new_n577), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G283), .B2(new_n852), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n268), .B1(new_n847), .B2(G107), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n601), .C2(new_n1037), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1106), .A2(KEYINPUT115), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(KEYINPUT115), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n268), .B1(new_n794), .B2(new_n402), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n800), .A2(new_n202), .B1(new_n796), .B2(new_n329), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G68), .C2(new_n852), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n816), .A2(G143), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n810), .A2(new_n858), .B1(new_n808), .B2(new_n861), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n821), .A2(G77), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1107), .A2(new_n1108), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1096), .B1(new_n1117), .B2(new_n787), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n786), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n983), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1092), .A2(new_n1093), .A3(new_n1120), .ZN(G390));
  OAI211_X1 g0921(.A(new_n361), .B(new_n705), .C1(new_n733), .C2(new_n737), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n869), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n898), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n926), .A2(new_n948), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n764), .A2(new_n898), .A3(new_n872), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1123), .B1(new_n875), .B2(new_n876), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n948), .B1(new_n1132), .B2(new_n898), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n947), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1130), .B(new_n1131), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n949), .B1(new_n959), .B2(new_n960), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n947), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n906), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n440), .B1(new_n930), .B2(new_n931), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n941), .B1(new_n1141), .B2(G330), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n872), .C1(new_n904), .C2(new_n905), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT117), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n960), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1143), .B2(new_n960), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1122), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1126), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1131), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n764), .A2(new_n872), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n960), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n959), .B1(new_n1139), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1142), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT118), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n440), .A2(new_n740), .ZN(new_n1156));
  INV_X1    g0956(.A(G330), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n696), .C1(new_n938), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1143), .A2(new_n960), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1143), .A2(new_n1144), .A3(new_n960), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1131), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1152), .B1(new_n906), .B2(new_n1157), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1132), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1158), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(G330), .A3(new_n1138), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT118), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1135), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1155), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n727), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1140), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n947), .A2(new_n782), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n841), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n771), .B1(new_n1176), .B2(new_n364), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n851), .B1(G283), .B2(new_n811), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n515), .B2(new_n808), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n268), .B(new_n1179), .C1(G87), .C2(new_n852), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n800), .A2(new_n345), .B1(new_n796), .B2(new_n443), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT120), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G294), .A2(new_n816), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1115), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n268), .B1(new_n794), .B2(new_n202), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n816), .B2(G125), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT119), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n852), .A2(new_n1064), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT53), .Z(new_n1190));
  NAND2_X1  g0990(.A1(new_n821), .A2(G159), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G132), .A2(new_n844), .B1(new_n801), .B2(G137), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT54), .B(G143), .Z(new_n1193));
  AOI22_X1  g0993(.A1(new_n811), .A2(G128), .B1(new_n826), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1185), .B1(new_n1188), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1177), .B1(new_n1196), .B2(new_n787), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1174), .A2(new_n770), .B1(new_n1175), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1173), .A2(new_n1198), .ZN(G378));
  NAND2_X1  g0999(.A1(new_n1171), .A2(new_n1142), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n371), .A2(new_n702), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n400), .A2(new_n384), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1204), .B1(new_n400), .B2(new_n384), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1202), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1207), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n1205), .A3(new_n1201), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n937), .B2(G330), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1211), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1157), .B(new_n1213), .C1(new_n927), .C2(new_n936), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n950), .B1(new_n962), .B2(new_n961), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT125), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n964), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n937), .A2(G330), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1213), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT125), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n937), .A2(G330), .A3(new_n1211), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1216), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1218), .A2(new_n1219), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1200), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1158), .B1(new_n1155), .B2(new_n1170), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1216), .A2(KEYINPUT124), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1215), .B(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1227), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n726), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n840), .B1(new_n841), .B2(new_n202), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n801), .A2(G97), .B1(new_n826), .B2(new_n505), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1234), .A2(KEYINPUT121), .B1(new_n855), .B2(new_n791), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n810), .A2(new_n515), .B1(new_n794), .B2(new_n416), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G107), .B2(new_n844), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G41), .B(new_n268), .C1(new_n852), .C2(G77), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1046), .A3(new_n1238), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1235), .B(new_n1239), .C1(KEYINPUT121), .C2(new_n1234), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT122), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT58), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(KEYINPUT58), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G33), .A2(G41), .ZN(new_n1244));
  AOI211_X1 g1044(.A(G50), .B(new_n1244), .C1(new_n342), .C2(new_n470), .ZN(new_n1245));
  INV_X1    g1045(.A(G128), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n808), .A2(new_n1246), .B1(new_n796), .B2(new_n860), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G125), .B2(new_n811), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G132), .A2(new_n801), .B1(new_n852), .B2(new_n1193), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n858), .C2(new_n1037), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n816), .A2(G124), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n1244), .C1(new_n861), .C2(new_n794), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1250), .B2(KEYINPUT59), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1245), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1242), .A2(new_n1243), .A3(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1233), .B1(new_n843), .B2(new_n1256), .C1(new_n1211), .C2(new_n783), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT123), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1230), .B2(new_n769), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1232), .A2(new_n1261), .ZN(G375));
  NAND3_X1  g1062(.A1(new_n1163), .A2(new_n1165), .A3(new_n1158), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1154), .A2(new_n998), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1193), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1265), .A2(new_n800), .B1(new_n860), .B2(new_n808), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n810), .A2(new_n854), .B1(new_n796), .B2(new_n858), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n818), .A2(new_n861), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n268), .B1(new_n794), .B2(new_n416), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1270), .B1(new_n202), .B2(new_n1037), .C1(new_n1246), .C2(new_n855), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n818), .A2(new_n443), .B1(new_n796), .B2(new_n345), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n268), .B(new_n1272), .C1(G77), .C2(new_n847), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n816), .A2(G303), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n810), .A2(new_n577), .B1(new_n808), .B2(new_n791), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n606), .B2(new_n801), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1066), .A3(new_n1274), .A4(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n843), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n771), .B1(new_n1176), .B2(G68), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1278), .B(new_n1279), .C1(new_n960), .C2(new_n782), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n770), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1264), .A2(new_n1282), .ZN(G381));
  AOI21_X1  g1083(.A(new_n1227), .B1(new_n1171), .B2(new_n1142), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n727), .B1(new_n1284), .B2(new_n1225), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1260), .B1(new_n1285), .B2(new_n1231), .ZN(new_n1286));
  INV_X1    g1086(.A(G378), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1052), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1290), .B(G390), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1291));
  NOR4_X1   g1091(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(KEYINPUT126), .ZN(G407));
  INV_X1    g1094(.A(G213), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1289), .B2(new_n703), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G407), .A2(new_n1296), .ZN(G409));
  XNOR2_X1  g1097(.A(G393), .B(new_n838), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(G390), .ZN(new_n1300));
  INV_X1    g1100(.A(G390), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1024), .A2(new_n1052), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1301), .B1(new_n1024), .B2(new_n1052), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1304), .A2(new_n1291), .A3(new_n1298), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G375), .A2(G378), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1295), .A2(G343), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1224), .A2(new_n1219), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1222), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n770), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AND4_X1   g1111(.A1(new_n1173), .A2(new_n1198), .A3(new_n1311), .A4(new_n1257), .ZN(new_n1312));
  OR3_X1    g1112(.A1(new_n1228), .A2(new_n1230), .A3(new_n999), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1308), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1307), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT60), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1263), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1263), .A2(new_n1316), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n726), .A3(new_n1154), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1282), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1319), .A2(G384), .A3(new_n1282), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(G2897), .A3(new_n1308), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1308), .A2(G2897), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1322), .A2(new_n1323), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1173), .A2(new_n1198), .A3(new_n1311), .A4(new_n1257), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1228), .A2(new_n1230), .A3(new_n999), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n1331), .A2(new_n1332), .B1(new_n1295), .B2(G343), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(G375), .B2(G378), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1324), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1335), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1314), .B(new_n1335), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1306), .A2(new_n1330), .A3(new_n1336), .A4(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1337), .A2(new_n1341), .A3(KEYINPUT62), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT62), .B1(new_n1337), .B2(new_n1341), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT61), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1334), .B2(new_n1328), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1342), .A2(new_n1343), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1340), .B1(new_n1346), .B2(new_n1306), .ZN(G405));
  NAND2_X1  g1147(.A1(new_n1307), .A2(new_n1288), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1335), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1307), .A2(new_n1288), .A3(new_n1324), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(new_n1306), .ZN(G402));
endmodule


