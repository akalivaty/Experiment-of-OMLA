//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT2), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  OAI211_X1 g008(.A(KEYINPUT79), .B(KEYINPUT2), .C1(new_n204), .C2(new_n205), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n203), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n209), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT2), .B2(new_n202), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT74), .B(G197gat), .ZN(new_n216));
  INV_X1    g015(.A(G204gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT22), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT22), .ZN(new_n221));
  INV_X1    g020(.A(G211gat), .ZN(new_n222));
  INV_X1    g021(.A(G218gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n225), .A2(KEYINPUT76), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(new_n225), .B2(KEYINPUT76), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT29), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n215), .B1(new_n229), .B2(KEYINPUT3), .ZN(new_n230));
  INV_X1    g029(.A(G228gat), .ZN(new_n231));
  INV_X1    g030(.A(G233gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n228), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n225), .A2(KEYINPUT76), .A3(new_n226), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n234), .A2(new_n235), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n230), .A2(new_n233), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n243), .A3(new_n226), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT81), .B1(new_n218), .B2(new_n224), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n216), .A2(G204gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n216), .A2(G204gat), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n246), .A2(KEYINPUT81), .A3(new_n247), .A4(new_n224), .ZN(new_n248));
  INV_X1    g047(.A(new_n226), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n244), .B(new_n236), .C1(new_n245), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n214), .B1(new_n251), .B2(new_n238), .ZN(new_n252));
  OAI22_X1  g051(.A1(new_n252), .A2(new_n240), .B1(new_n231), .B2(new_n232), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n242), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G78gat), .B(G106gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT31), .ZN(new_n256));
  INV_X1    g055(.A(G50gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT82), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n260), .A3(new_n253), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G22gat), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n253), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n259), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n254), .A2(new_n258), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n262), .A2(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(KEYINPUT64), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n274), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n277));
  INV_X1    g076(.A(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(G176gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT24), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(KEYINPUT24), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n270), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n285), .A2(KEYINPUT24), .ZN(new_n292));
  AND2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n292), .B1(new_n295), .B2(KEYINPUT24), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT25), .B1(new_n296), .B2(KEYINPUT67), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n273), .A2(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(KEYINPUT67), .A3(new_n287), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT68), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n270), .B1(new_n288), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n299), .A4(new_n298), .ZN(new_n305));
  OAI211_X1 g104(.A(KEYINPUT66), .B(new_n270), .C1(new_n283), .C2(new_n288), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n291), .A2(new_n301), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n272), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT26), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(KEYINPUT26), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n282), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT28), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT28), .B1(new_n312), .B2(new_n313), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n311), .B(new_n285), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT72), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n321), .A2(G113gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT70), .B(G113gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G120gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327));
  OR2_X1    g126(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT71), .B1(new_n330), .B2(new_n322), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n320), .A2(new_n326), .A3(new_n327), .A4(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(G127gat), .A2(G134gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT69), .B(G127gat), .Z(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  OAI221_X1 g135(.A(new_n333), .B1(new_n334), .B2(KEYINPUT1), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n307), .A2(new_n337), .A3(new_n332), .A4(new_n317), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT34), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n341), .A2(KEYINPUT34), .A3(new_n342), .ZN(new_n346));
  OAI211_X1 g145(.A(KEYINPUT32), .B(new_n343), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n341), .A2(new_n342), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT34), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(KEYINPUT32), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G71gat), .B(G99gat), .Z(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT73), .ZN(new_n356));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n347), .A2(new_n352), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n350), .A2(new_n344), .A3(new_n351), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n351), .B1(new_n350), .B2(new_n344), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n269), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n214), .A3(new_n337), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT4), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n332), .A2(new_n214), .A3(new_n369), .A4(new_n337), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n338), .B(new_n239), .C1(new_n375), .C2(new_n214), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n371), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n367), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n214), .B1(new_n332), .B2(new_n337), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n373), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n376), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n373), .A2(KEYINPUT5), .ZN(new_n383));
  OAI22_X1  g182(.A1(new_n377), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(G85gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391));
  OAI221_X1 g190(.A(new_n388), .B1(new_n382), .B2(new_n383), .C1(new_n377), .C2(new_n381), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT84), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n390), .A2(new_n396), .A3(new_n392), .A4(new_n391), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n318), .A2(KEYINPUT77), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n307), .A2(new_n401), .A3(new_n317), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n236), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n234), .A2(new_n235), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n318), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n318), .A2(KEYINPUT78), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n307), .A2(new_n401), .A3(new_n317), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n401), .B1(new_n307), .B2(new_n317), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n318), .A2(new_n236), .A3(new_n404), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n406), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  INV_X1    g220(.A(G64gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n399), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n417), .A2(new_n406), .A3(new_n418), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n403), .A2(new_n404), .B1(new_n411), .B2(new_n412), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n407), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n399), .A3(new_n430), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n366), .A2(new_n398), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n393), .A2(new_n395), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n414), .A2(new_n419), .A3(new_n430), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n414), .B2(new_n419), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n438), .A2(new_n439), .A3(new_n399), .ZN(new_n440));
  INV_X1    g239(.A(new_n433), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n365), .A2(KEYINPUT87), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n269), .A2(new_n444), .A3(new_n361), .A4(new_n364), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT35), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n436), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n265), .A2(new_n268), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n362), .A2(new_n363), .A3(new_n359), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n360), .B1(new_n347), .B2(new_n352), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n364), .A2(KEYINPUT36), .A3(new_n361), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n442), .A2(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n405), .A2(new_n406), .A3(new_n413), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n417), .A2(new_n407), .A3(new_n418), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT37), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n456), .B(new_n425), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n414), .A2(new_n461), .A3(new_n419), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n431), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT85), .B(new_n425), .C1(new_n429), .C2(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n414), .B2(new_n419), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(new_n430), .ZN(new_n467));
  INV_X1    g266(.A(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n398), .B(new_n463), .C1(new_n469), .C2(KEYINPUT38), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n382), .A2(new_n373), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT39), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(new_n389), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n378), .A2(new_n379), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n471), .B(KEYINPUT39), .C1(new_n373), .C2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n432), .A2(new_n390), .A3(new_n478), .A4(new_n433), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n473), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n269), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n455), .B1(new_n470), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n448), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n485));
  INV_X1    g284(.A(G29gat), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n488), .A2(new_n489), .B1(G29gat), .B2(G36gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(KEYINPUT15), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  XOR2_X1   g293(.A(G15gat), .B(G22gat), .Z(new_n495));
  INV_X1    g294(.A(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT16), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(G1gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n503), .A3(G8gat), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n497), .B(new_n502), .C1(new_n498), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n494), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT17), .B1(new_n494), .B2(KEYINPUT88), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n484), .B(new_n508), .C1(new_n513), .C2(new_n507), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT11), .B(G169gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G197gat), .ZN(new_n520));
  XOR2_X1   g319(.A(G113gat), .B(G141gat), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT12), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n508), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n509), .B(new_n510), .ZN(new_n527));
  INV_X1    g326(.A(new_n507), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT18), .A3(new_n484), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n494), .B(new_n507), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n484), .B(KEYINPUT13), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n530), .A2(new_n516), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n516), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(new_n518), .A3(new_n524), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n483), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT91), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n483), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  OR2_X1    g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G57gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(G64gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT92), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n422), .A2(G57gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT9), .B1(new_n552), .B2(new_n550), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n545), .A3(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n507), .B1(new_n557), .B2(KEYINPUT21), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G183gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G127gat), .B(G155gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT94), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n222), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n562), .A2(new_n565), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n566), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n566), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT95), .B(KEYINPUT97), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT96), .B(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n424), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n584), .A2(new_n585), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n591));
  INV_X1    g390(.A(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n494), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n590), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n581), .B(new_n594), .C1(new_n513), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(G134gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n527), .A2(new_n595), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(new_n336), .A3(new_n581), .A4(new_n594), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n580), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n205), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(new_n600), .A3(new_n580), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  INV_X1    g406(.A(new_n605), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(new_n601), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n544), .B1(new_n575), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(KEYINPUT98), .A3(new_n574), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n593), .A2(KEYINPUT100), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n557), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n595), .B2(new_n556), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n595), .A2(new_n620), .A3(new_n556), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n618), .B(new_n619), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n557), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n279), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n217), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n543), .A2(new_n614), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n437), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n496), .ZN(G1324gat));
  NOR2_X1   g440(.A1(new_n639), .A2(new_n434), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n501), .A2(new_n505), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n501), .A2(new_n505), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(G8gat), .B1(new_n639), .B2(new_n434), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n642), .A2(KEYINPUT42), .A3(new_n644), .A4(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(G1325gat));
  INV_X1    g450(.A(new_n639), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n453), .A2(new_n454), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(G15gat), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G15gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n451), .A2(new_n452), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n639), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n655), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(G1326gat));
  NOR2_X1   g463(.A1(new_n639), .A2(new_n269), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT43), .B(G22gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  INV_X1    g466(.A(new_n638), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n574), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n541), .B1(new_n483), .B2(new_n538), .ZN(new_n670));
  INV_X1    g469(.A(new_n538), .ZN(new_n671));
  AOI211_X1 g470(.A(KEYINPUT91), .B(new_n671), .C1(new_n448), .C2(new_n482), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n610), .B(new_n669), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n437), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n486), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n482), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(KEYINPUT102), .B(new_n455), .C1(new_n470), .C2(new_n481), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n448), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n681), .B2(new_n610), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  AOI211_X1 g482(.A(new_n683), .B(new_n612), .C1(new_n448), .C2(new_n482), .ZN(new_n684));
  INV_X1    g483(.A(new_n669), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n682), .A2(new_n684), .A3(new_n671), .A4(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(new_n675), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n486), .B2(new_n687), .ZN(G1328gat));
  NOR3_X1   g487(.A1(new_n673), .A2(G36gat), .A3(new_n434), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  INV_X1    g489(.A(new_n434), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n686), .A2(KEYINPUT103), .A3(new_n691), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(G36gat), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n690), .A2(new_n696), .ZN(G1329gat));
  NAND3_X1  g496(.A1(new_n686), .A2(G43gat), .A3(new_n654), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT47), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n673), .B2(new_n658), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n699), .A2(KEYINPUT47), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1330gat));
  AOI21_X1  g504(.A(new_n257), .B1(new_n686), .B2(new_n449), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n269), .A2(G50gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT105), .Z(new_n709));
  NOR2_X1   g508(.A1(new_n673), .A2(new_n709), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n706), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1331gat));
  NAND3_X1  g512(.A1(new_n614), .A2(new_n668), .A3(new_n671), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n681), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n437), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n549), .ZN(G1332gat));
  INV_X1    g517(.A(new_n716), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n434), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n719), .B(new_n720), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT49), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n722), .B(new_n422), .C1(new_n716), .C2(new_n434), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n721), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n719), .A2(G71gat), .A3(new_n654), .ZN(new_n728));
  INV_X1    g527(.A(G71gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n716), .B2(new_n658), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n719), .A2(new_n449), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n681), .A2(new_n610), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n684), .B1(new_n736), .B2(new_n683), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n574), .A2(new_n538), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n668), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n735), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NOR4_X1   g540(.A1(new_n682), .A2(new_n684), .A3(KEYINPUT109), .A4(new_n739), .ZN(new_n742));
  OAI211_X1 g541(.A(G85gat), .B(new_n675), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n738), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT51), .B1(new_n736), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n681), .A2(new_n746), .A3(new_n610), .A4(new_n738), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n745), .A2(new_n675), .A3(new_n668), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n587), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1336gat));
  NAND4_X1  g553(.A1(new_n745), .A2(new_n668), .A3(new_n691), .A4(new_n747), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(G92gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n691), .B1(new_n741), .B2(new_n742), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G92gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n737), .A2(new_n740), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n434), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n737), .A2(KEYINPUT111), .A3(new_n691), .A4(new_n740), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n762), .A2(G92gat), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n759), .B1(new_n755), .B2(G92gat), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n758), .A2(new_n759), .B1(new_n764), .B2(new_n765), .ZN(G1337gat));
  NOR2_X1   g565(.A1(new_n741), .A2(new_n742), .ZN(new_n767));
  OAI21_X1  g566(.A(G99gat), .B1(new_n767), .B2(new_n653), .ZN(new_n768));
  INV_X1    g567(.A(G99gat), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n745), .A2(new_n769), .A3(new_n668), .A4(new_n747), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n658), .B2(new_n770), .ZN(G1338gat));
  OAI211_X1 g570(.A(KEYINPUT53), .B(G106gat), .C1(new_n767), .C2(new_n269), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n269), .A2(G106gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n745), .A2(new_n668), .A3(new_n747), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT112), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G106gat), .B1(new_n761), .B2(new_n269), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n774), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n772), .A2(new_n777), .B1(new_n780), .B2(new_n775), .ZN(G1339gat));
  NAND3_X1  g580(.A1(new_n623), .A2(new_n629), .A3(new_n624), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n623), .A2(KEYINPUT113), .A3(new_n629), .A4(new_n624), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n784), .A2(new_n627), .A3(KEYINPUT54), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n629), .B1(new_n623), .B2(new_n624), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n636), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n637), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n786), .A2(new_n789), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(KEYINPUT114), .A3(new_n637), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n793), .A2(new_n538), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n529), .A2(new_n484), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n531), .A2(new_n532), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n522), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n536), .B2(new_n524), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n802), .A2(new_n638), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n610), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n610), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n801), .B(KEYINPUT115), .C1(new_n536), .C2(new_n524), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n796), .A3(new_n797), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n575), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n611), .A2(new_n613), .A3(new_n638), .A4(new_n671), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT116), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n366), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n691), .A2(new_n437), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n671), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n443), .A2(new_n445), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n817), .A2(new_n675), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n434), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n538), .A2(new_n323), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n820), .B2(new_n638), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n321), .A3(new_n434), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n638), .ZN(G1341gat));
  NOR3_X1   g630(.A1(new_n820), .A2(new_n335), .A3(new_n575), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n825), .A2(new_n574), .A3(new_n434), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n335), .ZN(G1342gat));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n612), .A2(G134gat), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n825), .A2(new_n835), .A3(new_n434), .A4(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n817), .A2(new_n822), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n824), .A3(new_n675), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n434), .A3(new_n840), .A4(new_n836), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n820), .B2(new_n612), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  INV_X1    g645(.A(new_n791), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n786), .B2(new_n789), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n795), .B1(new_n794), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n538), .B(new_n847), .C1(new_n848), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n610), .B1(new_n851), .B2(new_n803), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n575), .B1(new_n852), .B2(new_n810), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n846), .B(new_n269), .C1(new_n853), .C2(new_n812), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n815), .A2(new_n449), .A3(new_n816), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(G141gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n819), .A2(new_n653), .ZN(new_n860));
  NOR4_X1   g659(.A1(new_n858), .A2(new_n859), .A3(new_n671), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n855), .A2(new_n860), .ZN(new_n862));
  AOI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n538), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n845), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n845), .B(new_n866), .C1(new_n861), .C2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  NAND4_X1  g667(.A1(new_n815), .A2(new_n449), .A3(new_n816), .A4(new_n856), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n853), .A2(new_n812), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n846), .B1(new_n870), .B2(new_n269), .ZN(new_n871));
  AOI211_X1 g670(.A(new_n638), .B(new_n860), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT59), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  INV_X1    g674(.A(new_n854), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n815), .A2(new_n449), .A3(new_n816), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n856), .ZN(new_n878));
  INV_X1    g677(.A(new_n860), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n880), .B2(new_n638), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n874), .B1(new_n881), .B2(new_n873), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n862), .A2(new_n873), .A3(new_n668), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n574), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n204), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n574), .A2(G155gat), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT121), .Z(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n880), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(G1346gat));
  NOR3_X1   g690(.A1(new_n880), .A2(new_n205), .A3(new_n612), .ZN(new_n892));
  AOI21_X1  g691(.A(G162gat), .B1(new_n862), .B2(new_n610), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n434), .A2(new_n675), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n838), .A2(new_n278), .A3(new_n538), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n817), .A2(new_n366), .A3(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n671), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT123), .ZN(G1348gat));
  NOR3_X1   g699(.A1(new_n897), .A2(new_n279), .A3(new_n638), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n838), .A2(new_n668), .A3(new_n895), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n279), .B2(new_n902), .ZN(G1349gat));
  NAND4_X1  g702(.A1(new_n838), .A2(new_n574), .A3(new_n312), .A4(new_n895), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n897), .B2(new_n575), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT124), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n906), .B(new_n908), .ZN(G1350gat));
  NAND4_X1  g708(.A1(new_n838), .A2(new_n313), .A3(new_n610), .A4(new_n895), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n818), .A2(new_n610), .A3(new_n895), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(G190gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n911), .B2(G190gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n869), .A2(new_n871), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n653), .A2(new_n895), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n671), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n855), .A2(new_n918), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n538), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1352gat));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n877), .A2(new_n217), .A3(new_n668), .A4(new_n919), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(KEYINPUT62), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n855), .A2(new_n918), .A3(G204gat), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n929), .A2(KEYINPUT125), .A3(new_n930), .A4(new_n668), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n638), .B(new_n918), .C1(new_n869), .C2(new_n871), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n217), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n668), .A3(new_n919), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n937), .A2(G204gat), .B1(new_n927), .B2(KEYINPUT62), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n928), .A4(new_n931), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n940), .ZN(G1353gat));
  OAI21_X1  g740(.A(G211gat), .B1(new_n920), .B2(new_n575), .ZN(new_n942));
  NAND2_X1  g741(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n943));
  OR2_X1    g742(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n922), .A2(new_n222), .A3(new_n574), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n945), .B(new_n946), .C1(new_n942), .C2(new_n944), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n920), .B2(new_n612), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n922), .A2(new_n223), .A3(new_n610), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1355gat));
endmodule


