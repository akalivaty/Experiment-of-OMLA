//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n452, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G234));
  INV_X1    g026(.A(G2106), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  OAI22_X1  g035(.A1(new_n456), .A2(new_n452), .B1(new_n449), .B2(new_n457), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT70), .B1(new_n464), .B2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(new_n473), .A2(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT71), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n485), .A2(KEYINPUT71), .A3(new_n486), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n465), .A3(new_n467), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n473), .A2(G138), .A3(new_n474), .A4(new_n475), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n475), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n499), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(new_n513), .A3(G62), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n505), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n517), .A2(new_n523), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n525), .A2(new_n531), .ZN(G168));
  INV_X1    g107(.A(new_n517), .ZN(new_n533));
  INV_X1    g108(.A(new_n519), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G90), .B1(G52), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n507), .A2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(KEYINPUT74), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n534), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OAI221_X1 g121(.A(new_n544), .B1(new_n545), .B2(new_n517), .C1(new_n546), .C2(new_n505), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT75), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND4_X1  g129(.A1(new_n516), .A2(KEYINPUT76), .A3(G53), .A4(G543), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n505), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n533), .A2(KEYINPUT77), .A3(G91), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n517), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n556), .A2(new_n558), .A3(new_n559), .A4(new_n562), .ZN(G299));
  XNOR2_X1  g138(.A(new_n542), .B(KEYINPUT78), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n533), .A2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n534), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  AOI22_X1  g145(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n505), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n517), .A2(new_n573), .B1(new_n519), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n572), .A2(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(G72), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G60), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n537), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(G651), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n533), .A2(G85), .B1(G47), .B2(new_n534), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G290));
  AND3_X1   g162(.A1(new_n510), .A2(G92), .A3(new_n516), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n537), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(G54), .A2(new_n534), .B1(new_n592), .B2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G301), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n595), .ZN(G284));
  XNOR2_X1  g173(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g174(.A1(G299), .A2(new_n595), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n595), .B2(G168), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(new_n595), .B2(G168), .ZN(G280));
  INV_X1    g177(.A(new_n594), .ZN(new_n603));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n483), .A2(G135), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT82), .ZN(new_n611));
  INV_X1    g186(.A(new_n485), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n474), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT83), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT12), .Z(new_n620));
  XOR2_X1   g195(.A(KEYINPUT13), .B(G2100), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(G401));
  XNOR2_X1  g214(.A(G2072), .B(G2078), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT85), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2096), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n642), .A2(new_n643), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n650), .B2(new_n644), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n648), .B(new_n651), .Z(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n657), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  OAI221_X1 g237(.A(new_n658), .B1(new_n655), .B2(new_n659), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G1991), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G16), .A2(G23), .ZN(new_n672));
  INV_X1    g247(.A(G288), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n673), .B2(G16), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT33), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G22), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G166), .B2(new_n677), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G1971), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(G1971), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(G6), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n572), .A2(new_n575), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n677), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n676), .A2(new_n680), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT34), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n677), .A2(G24), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n690), .B(new_n691), .C1(G290), .C2(G16), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G1986), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n612), .A2(KEYINPUT88), .A3(G119), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G131), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n697));
  INV_X1    g272(.A(G119), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n485), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n695), .A2(new_n696), .A3(new_n699), .A4(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT35), .B(G1991), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  OR2_X1    g280(.A1(new_n693), .A2(G1986), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n688), .A2(new_n694), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT36), .ZN(new_n708));
  NAND2_X1  g283(.A1(G171), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G5), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT95), .ZN(new_n713));
  NAND2_X1  g288(.A1(G168), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G21), .ZN(new_n715));
  INV_X1    g290(.A(G1966), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT94), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(G28), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(G28), .ZN(new_n722));
  AND2_X1   g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  NOR2_X1   g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n720), .A2(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n715), .B2(new_n716), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n713), .B(new_n727), .C1(new_n721), .C2(new_n617), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT96), .Z(new_n729));
  AND2_X1   g304(.A1(new_n710), .A2(new_n711), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(KEYINPUT24), .B2(G34), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(KEYINPUT24), .B2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n479), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2084), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n677), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n548), .B2(new_n677), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n736), .B2(G1341), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n730), .B(new_n737), .C1(G1341), .C2(new_n736), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n483), .A2(G141), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n612), .A2(G129), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(G105), .B2(new_n477), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n739), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n749), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n677), .A2(G4), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n603), .B2(new_n677), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1348), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n477), .A2(G103), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n465), .A2(new_n467), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n759), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  INV_X1    g335(.A(G139), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n758), .B1(new_n474), .B2(new_n760), .C1(new_n482), .C2(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G33), .B(new_n762), .S(G29), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2072), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n752), .A2(new_n755), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G299), .A2(G16), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n677), .A2(G20), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(G162), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G29), .B2(G35), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2090), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n738), .A2(new_n765), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n721), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n782));
  INV_X1    g357(.A(G140), .ZN(new_n783));
  INV_X1    g358(.A(G128), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n782), .B1(new_n482), .B2(new_n783), .C1(new_n784), .C2(new_n485), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n787), .A2(KEYINPUT91), .A3(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT91), .B1(new_n787), .B2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n780), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  NOR2_X1   g366(.A1(G27), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT97), .B(G2078), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n774), .B2(new_n776), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n778), .A2(new_n791), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n708), .A2(new_n729), .A3(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  AOI22_X1  g375(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n505), .ZN(new_n802));
  INV_X1    g377(.A(G93), .ZN(new_n803));
  INV_X1    g378(.A(G55), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n517), .A2(new_n803), .B1(new_n519), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G860), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT37), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n547), .A2(new_n806), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n806), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n548), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n603), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(G860), .B1(new_n818), .B2(KEYINPUT39), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n819), .A2(new_n820), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n809), .B1(new_n823), .B2(new_n824), .ZN(G145));
  INV_X1    g400(.A(G164), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n787), .B(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n747), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n747), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n762), .B(KEYINPUT102), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n828), .A2(KEYINPUT102), .A3(new_n762), .A4(new_n829), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n702), .B(new_n620), .ZN(new_n834));
  OR2_X1    g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G118), .C2(new_n474), .ZN(new_n836));
  INV_X1    g411(.A(G142), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n482), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G130), .B2(new_n612), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n834), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT103), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(KEYINPUT103), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n832), .A2(new_n833), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n617), .B(new_n479), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n832), .A2(new_n833), .A3(new_n840), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  AND4_X1   g424(.A1(new_n833), .A2(new_n832), .A3(new_n842), .A4(new_n841), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(new_n843), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n848), .B(new_n849), .C1(new_n851), .C2(new_n846), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g428(.A1(new_n603), .A2(G299), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT105), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n603), .A2(G299), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(KEYINPUT105), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n855), .A2(KEYINPUT41), .A3(new_n856), .A4(new_n857), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(KEYINPUT106), .A3(new_n861), .ZN(new_n862));
  OR3_X1    g437(.A1(new_n858), .A2(KEYINPUT106), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n606), .B(KEYINPUT104), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n813), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n858), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT42), .ZN(new_n869));
  XNOR2_X1  g444(.A(G290), .B(G288), .ZN(new_n870));
  XNOR2_X1  g445(.A(G166), .B(new_n683), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n870), .B(new_n871), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(KEYINPUT107), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(KEYINPUT42), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n869), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n869), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(G868), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n812), .A2(new_n595), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(G295));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n879), .ZN(G331));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n882));
  INV_X1    g457(.A(new_n813), .ZN(new_n883));
  NAND2_X1  g458(.A1(G301), .A2(G168), .ZN(new_n884));
  NAND2_X1  g459(.A1(G171), .A2(G286), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT108), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n813), .A2(new_n884), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n890), .B2(KEYINPUT108), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n858), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n860), .A2(KEYINPUT109), .A3(new_n861), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n858), .A2(KEYINPUT109), .A3(new_n859), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n890), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n873), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n888), .A2(new_n858), .A3(new_n889), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n873), .B(new_n898), .C1(new_n864), .C2(new_n891), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n897), .A2(new_n899), .A3(new_n900), .A4(new_n849), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n849), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT110), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n882), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n898), .B1(new_n864), .B2(new_n891), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n905), .A2(new_n872), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(new_n902), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT44), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n897), .A2(new_n882), .A3(new_n849), .A4(new_n899), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n907), .B2(new_n882), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(G397));
  INV_X1    g489(.A(KEYINPUT127), .ZN(new_n915));
  INV_X1    g490(.A(G1384), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n499), .B2(new_n503), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n471), .A2(G40), .A3(new_n476), .A4(new_n478), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(KEYINPUT45), .B(new_n916), .C1(new_n499), .C2(new_n503), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(KEYINPUT50), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT50), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(new_n916), .C1(new_n499), .C2(new_n503), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n926), .A3(new_n921), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n923), .A2(G1966), .B1(G2084), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(G8), .ZN(new_n929));
  INV_X1    g504(.A(G8), .ZN(new_n930));
  NOR2_X1   g505(.A1(G168), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(KEYINPUT51), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT51), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n935), .B(G8), .C1(new_n928), .C2(G286), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n937), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT126), .B1(new_n937), .B2(KEYINPUT62), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n922), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n919), .ZN(new_n943));
  INV_X1    g518(.A(G2078), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n917), .A2(new_n941), .A3(new_n918), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n921), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT53), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n927), .A2(new_n711), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(G2078), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n919), .A2(new_n921), .A3(new_n922), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n597), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n937), .B2(KEYINPUT62), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n943), .A2(new_n921), .A3(new_n945), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(G1971), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n927), .A2(G2090), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n957), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n920), .B1(new_n942), .B2(new_n919), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n945), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT114), .B1(new_n965), .B2(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G166), .B2(new_n930), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT55), .B(G8), .C1(new_n515), .C2(new_n521), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(KEYINPUT115), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n962), .A2(new_n966), .A3(G8), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(G8), .B1(new_n965), .B2(new_n960), .ZN(new_n976));
  INV_X1    g551(.A(new_n970), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n979));
  NOR2_X1   g554(.A1(G305), .A2(G1981), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n683), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT49), .ZN(new_n984));
  INV_X1    g559(.A(new_n917), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n930), .B1(new_n985), .B2(new_n921), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n979), .B(new_n987), .C1(new_n980), .C2(new_n982), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n673), .A2(G1976), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT52), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n989), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n975), .A2(new_n978), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT123), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n975), .A2(KEYINPUT123), .A3(new_n996), .A4(new_n978), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n955), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT125), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n940), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT125), .B(new_n955), .C1(new_n999), .C2(new_n1000), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n915), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n999), .A2(new_n1000), .ZN(new_n1006));
  INV_X1    g581(.A(new_n955), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT125), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(KEYINPUT127), .A3(new_n1010), .A4(new_n940), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT63), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n928), .A2(G8), .A3(G168), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n997), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n962), .A2(new_n966), .A3(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n977), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1013), .A2(new_n1012), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(new_n975), .A3(new_n996), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n975), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n989), .A2(new_n991), .A3(new_n673), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(G1981), .B2(G305), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1020), .A2(new_n996), .B1(new_n1022), .B2(new_n986), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n999), .A2(new_n1000), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1025));
  XNOR2_X1  g600(.A(G299), .B(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n943), .A2(new_n921), .A3(new_n945), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1956), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n927), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n917), .A2(G2067), .A3(new_n920), .ZN(new_n1032));
  INV_X1    g607(.A(G1348), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n927), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT118), .B1(new_n1034), .B2(new_n594), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n920), .B1(new_n917), .B2(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1348), .B1(new_n1037), .B2(new_n926), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1036), .B(new_n603), .C1(new_n1038), .C2(new_n1032), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1028), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1031), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1996), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n1043), .A2(new_n943), .A3(new_n921), .A4(new_n945), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n917), .B2(new_n920), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n548), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT59), .B(new_n548), .C1(new_n1044), .C2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1041), .B1(KEYINPUT120), .B2(KEYINPUT61), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1034), .A2(KEYINPUT60), .A3(new_n594), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1056));
  AND2_X1   g631(.A1(new_n1034), .A2(KEYINPUT60), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n603), .B1(new_n1034), .B2(KEYINPUT60), .ZN(new_n1058));
  OAI221_X1 g633(.A(new_n1055), .B1(new_n1041), .B2(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1042), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n950), .B1(new_n920), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1063), .B2(new_n920), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n919), .A2(new_n922), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n949), .A2(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n927), .A2(KEYINPUT121), .A3(new_n711), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n948), .A3(G301), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n953), .A2(new_n1061), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n948), .A3(new_n1068), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n949), .A2(new_n951), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n947), .B2(new_n946), .ZN(new_n1073));
  AOI22_X1  g648(.A1(G171), .A2(new_n1071), .B1(new_n1073), .B2(G301), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1070), .B1(new_n1074), .B2(new_n1061), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1060), .A2(new_n1075), .A3(new_n937), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1019), .B(new_n1023), .C1(new_n1024), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1006), .A2(new_n937), .A3(new_n1060), .A4(new_n1075), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(KEYINPUT124), .A3(new_n1019), .A4(new_n1023), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1005), .A2(new_n1011), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n919), .A2(new_n920), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1043), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n747), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(KEYINPUT111), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(KEYINPUT111), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n787), .B(G2067), .Z(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1043), .B2(new_n748), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1087), .B(new_n1088), .C1(new_n1090), .C2(new_n1083), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n702), .A2(new_n704), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n702), .A2(new_n704), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G290), .B(G1986), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1083), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1082), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1083), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n787), .A2(G2067), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1089), .A2(new_n748), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT46), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1103), .A2(new_n1083), .B1(new_n1104), .B2(new_n1084), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1104), .B2(new_n1084), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT47), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1095), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1099), .A2(G290), .A3(G1986), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT48), .Z(new_n1111));
  AOI211_X1 g686(.A(new_n1102), .B(new_n1108), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1098), .A2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g688(.A(G319), .ZN(new_n1115));
  NOR3_X1   g689(.A1(G401), .A2(new_n1115), .A3(G227), .ZN(new_n1116));
  NAND4_X1  g690(.A1(new_n911), .A2(new_n852), .A3(new_n670), .A4(new_n1116), .ZN(G225));
  INV_X1    g691(.A(G225), .ZN(G308));
endmodule


