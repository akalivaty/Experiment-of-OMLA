//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(G472), .B2(G902), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT32), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT31), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AND4_X1   g019(.A1(new_n198), .A2(new_n203), .A3(new_n205), .A4(new_n200), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(G143), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(KEYINPUT64), .A3(G146), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n208), .A2(new_n209), .B1(G143), .B2(new_n202), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n200), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n201), .A2(new_n206), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G137), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT66), .B(new_n215), .C1(new_n216), .C2(G137), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G134), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT11), .A4(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n221), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n220), .ZN(new_n230));
  INV_X1    g044(.A(G131), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n226), .A4(new_n227), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n214), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT2), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n199), .A2(new_n251), .A3(G128), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n210), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n216), .A2(G137), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n223), .A2(G134), .ZN(new_n257));
  OAI21_X1  g071(.A(G131), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n232), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n233), .A2(new_n250), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT30), .B1(new_n233), .B2(new_n259), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n199), .A2(new_n200), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n199), .A2(new_n198), .A3(new_n200), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n208), .A2(new_n209), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n203), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n263), .A2(new_n264), .B1(new_n266), .B2(new_n212), .ZN(new_n267));
  INV_X1    g081(.A(new_n232), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n226), .A2(new_n227), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n231), .B1(new_n269), .B2(new_n230), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n232), .A2(new_n255), .A3(new_n258), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n261), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n260), .B1(new_n275), .B2(new_n248), .ZN(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n278), .B(KEYINPUT27), .Z(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n197), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n261), .A2(new_n274), .B1(new_n240), .B2(new_n247), .ZN(new_n284));
  NOR4_X1   g098(.A1(new_n284), .A2(KEYINPUT31), .A3(new_n260), .A4(new_n281), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n271), .A2(new_n273), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n250), .B1(new_n287), .B2(KEYINPUT69), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n233), .A2(new_n259), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT28), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n248), .ZN(new_n294));
  INV_X1    g108(.A(new_n250), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n281), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n196), .B1(new_n286), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n275), .A2(new_n248), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n296), .A3(new_n282), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT31), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n276), .A2(new_n197), .A3(new_n282), .ZN(new_n303));
  AND4_X1   g117(.A1(new_n196), .A2(new_n302), .A3(new_n298), .A4(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n195), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n192), .B1(new_n299), .B2(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n194), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n302), .A2(new_n298), .A3(new_n303), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT70), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n302), .A2(new_n298), .A3(new_n196), .A4(new_n303), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n195), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n282), .B1(new_n292), .B2(new_n297), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n276), .A2(new_n281), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n287), .A2(new_n250), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n296), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n292), .B1(KEYINPUT28), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n281), .A2(new_n318), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n187), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n307), .A2(new_n309), .A3(new_n314), .A4(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G214), .B1(G237), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(G952), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G953), .ZN(new_n330));
  INV_X1    g144(.A(G234), .ZN(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G953), .ZN(new_n335));
  AOI211_X1 g149(.A(new_n188), .B(new_n335), .C1(G234), .C2(G237), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT21), .B(G898), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n204), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n253), .A2(G143), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n339), .A2(new_n340), .A3(new_n216), .ZN(new_n341));
  XNOR2_X1  g155(.A(G116), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G107), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT13), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n340), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n339), .A2(new_n348), .ZN(new_n351));
  OAI21_X1  g165(.A(G134), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n243), .A2(KEYINPUT14), .A3(G122), .ZN(new_n354));
  OAI211_X1 g168(.A(G107), .B(new_n354), .C1(new_n343), .C2(KEYINPUT14), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n216), .B1(new_n339), .B2(new_n340), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n355), .B(new_n346), .C1(new_n341), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT9), .B(G234), .ZN(new_n359));
  INV_X1    g173(.A(G217), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n359), .A2(new_n360), .A3(G953), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n357), .A3(new_n361), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G478), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n365), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(G125), .A3(G140), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(KEYINPUT16), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(G125), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G146), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n202), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n332), .A2(new_n335), .A3(G214), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n204), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n277), .A2(G143), .A3(G214), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n231), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n231), .B1(new_n385), .B2(new_n386), .ZN(new_n389));
  OR3_X1    g203(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT17), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n379), .A2(KEYINPUT93), .A3(new_n380), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(KEYINPUT17), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n383), .A2(new_n390), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n386), .ZN(new_n394));
  AOI21_X1  g208(.A(G143), .B1(new_n277), .B2(G214), .ZN(new_n395));
  OAI211_X1 g209(.A(KEYINPUT18), .B(G131), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n371), .A2(G146), .A3(new_n373), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n370), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n375), .A2(new_n398), .A3(new_n202), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT18), .A2(G131), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n385), .A2(new_n386), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n396), .A2(KEYINPUT89), .A3(new_n402), .A4(new_n400), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G113), .B(G122), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT92), .B(G104), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n393), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n393), .B2(new_n407), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n188), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G475), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n371), .A2(KEYINPUT19), .A3(new_n373), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT19), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n375), .A2(new_n398), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT91), .B1(new_n419), .B2(G146), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n416), .A2(new_n421), .A3(new_n418), .A4(new_n202), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n389), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT90), .A3(new_n387), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n388), .B2(new_n389), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n423), .A2(new_n425), .A3(new_n427), .A4(new_n379), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n407), .ZN(new_n429));
  INV_X1    g243(.A(new_n410), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n393), .A2(new_n407), .A3(new_n410), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n415), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  AOI211_X1 g250(.A(KEYINPUT20), .B(new_n436), .C1(new_n431), .C2(new_n432), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n414), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n414), .B(KEYINPUT94), .C1(new_n435), .C2(new_n437), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n338), .B(new_n368), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT8), .ZN(new_n444));
  INV_X1    g258(.A(G101), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n345), .A2(G104), .ZN(new_n446));
  INV_X1    g260(.A(G104), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT3), .B1(new_n447), .B2(G107), .ZN(new_n450));
  AOI21_X1  g264(.A(G101), .B1(new_n447), .B2(G107), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT3), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n345), .A3(G104), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT80), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n450), .A2(new_n451), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n449), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n234), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n460), .A2(new_n461), .B1(new_n239), .B2(new_n238), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n458), .A2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n444), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n335), .A2(G224), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(KEYINPUT86), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(KEYINPUT86), .B2(new_n468), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n267), .A2(new_n370), .ZN(new_n471));
  INV_X1    g285(.A(new_n254), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n266), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n370), .A3(new_n252), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n470), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n474), .B(new_n466), .C1(new_n267), .C2(new_n370), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n478), .A2(new_n468), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n470), .C1(new_n471), .C2(new_n475), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n465), .A2(new_n477), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n458), .A2(new_n462), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n455), .A2(new_n457), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n450), .A2(new_n453), .A3(new_n448), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(G101), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(G101), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n248), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n443), .B(new_n483), .C1(new_n488), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT84), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n487), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n248), .A2(new_n490), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n494), .A2(new_n495), .B1(new_n458), .B2(new_n462), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n443), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n482), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n496), .B2(new_n443), .ZN(new_n504));
  INV_X1    g318(.A(new_n443), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n491), .B1(new_n484), .B2(new_n487), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n505), .B(new_n502), .C1(new_n506), .C2(new_n463), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n498), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n467), .B1(new_n471), .B2(new_n475), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(new_n478), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT85), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n515), .B(new_n512), .C1(new_n508), .C2(new_n509), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n500), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n518));
  OAI21_X1  g332(.A(G210), .B1(G237), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n520), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n519), .B(new_n500), .C1(new_n514), .C2(new_n516), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(KEYINPUT88), .A3(new_n523), .ZN(new_n524));
  AND4_X1   g338(.A1(new_n328), .A2(new_n442), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT24), .B(G110), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT74), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n241), .A2(G128), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n241), .A2(G128), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n531), .B(new_n535), .C1(new_n528), .C2(KEYINPUT23), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n536), .A2(G110), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n533), .B2(new_n537), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n399), .B(new_n379), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(G110), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n381), .B(new_n541), .C1(new_n527), .C2(new_n532), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT22), .B(G137), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n335), .A2(G221), .A3(G234), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n547), .B(new_n548), .Z(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n540), .B(new_n549), .C1(new_n544), .C2(new_n545), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G217), .B1(new_n331), .B2(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n188), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n554), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n561), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n551), .A2(new_n552), .A3(new_n563), .A4(new_n559), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n556), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(KEYINPUT79), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT79), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n567), .B(new_n556), .C1(new_n562), .C2(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n229), .A2(new_n232), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n252), .B1(new_n199), .B2(new_n254), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n458), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n458), .A2(new_n255), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n458), .A2(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n570), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n494), .A2(new_n267), .A3(new_n490), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n458), .A2(KEYINPUT10), .A3(new_n255), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G140), .ZN(new_n583));
  INV_X1    g397(.A(G227), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G953), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n575), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n570), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n587), .B1(new_n591), .B2(new_n582), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n569), .B(new_n188), .C1(new_n589), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n582), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n586), .B1(new_n575), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n582), .A2(KEYINPUT82), .A3(new_n587), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(G469), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(G469), .A2(G902), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n593), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G221), .B1(new_n359), .B2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n566), .A2(new_n568), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n327), .A2(new_n525), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n522), .A2(new_n608), .A3(new_n523), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n328), .B1(new_n523), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT96), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n338), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n440), .A2(new_n441), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  INV_X1    g428(.A(new_n364), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n361), .B1(new_n353), .B2(new_n357), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n614), .B(new_n366), .C1(new_n617), .C2(G902), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT98), .B1(new_n365), .B2(G478), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n358), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n617), .A2(KEYINPUT33), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(KEYINPUT33), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n615), .B2(new_n616), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n366), .A2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n620), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n621), .B1(new_n620), .B2(new_n628), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n328), .ZN(new_n634));
  INV_X1    g448(.A(new_n523), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(KEYINPUT95), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n522), .A2(new_n608), .A3(new_n523), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n611), .A2(new_n612), .A3(new_n633), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n193), .B1(new_n311), .B2(new_n312), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n313), .A2(new_n188), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(G472), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n605), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT100), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(new_n368), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n438), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n611), .A2(new_n612), .A3(new_n639), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n645), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  INV_X1    g470(.A(new_n604), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n562), .A2(new_n564), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n546), .B(new_n659), .Z(new_n660));
  OAI21_X1  g474(.A(new_n658), .B1(new_n555), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n525), .A2(new_n644), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n327), .A2(new_n663), .ZN(new_n668));
  INV_X1    g482(.A(new_n336), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n333), .B1(new_n669), .B2(G900), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n651), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n611), .A2(new_n639), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n667), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT72), .B1(new_n313), .B2(new_n195), .ZN(new_n674));
  INV_X1    g488(.A(new_n195), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n306), .B(new_n675), .C1(new_n311), .C2(new_n312), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n325), .B1(new_n308), .B2(new_n194), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n662), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n637), .B1(new_n636), .B2(new_n638), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(new_n682), .A3(KEYINPUT101), .A4(new_n671), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XNOR2_X1  g499(.A(new_n670), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n657), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n613), .A2(new_n650), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n688), .A2(new_n689), .A3(new_n634), .A4(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n276), .A2(new_n281), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n188), .B1(new_n321), .B2(new_n282), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n308), .A2(new_n194), .B1(G472), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n677), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n661), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n524), .A2(new_n521), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n692), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NAND2_X1  g517(.A1(new_n633), .A2(new_n670), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n611), .A2(new_n705), .A3(new_n639), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n668), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n202), .ZN(G48));
  NOR2_X1   g522(.A1(new_n566), .A2(new_n568), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n589), .A2(new_n592), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n593), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n603), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n327), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n640), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT41), .B(G113), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NOR2_X1   g533(.A1(new_n716), .A2(new_n652), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n243), .ZN(G18));
  AND2_X1   g535(.A1(new_n442), .A2(new_n661), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n307), .A2(new_n314), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n326), .B1(new_n642), .B2(KEYINPUT32), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n611), .A2(new_n639), .A3(new_n715), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n241), .ZN(G21));
  NAND3_X1  g542(.A1(new_n611), .A2(new_n639), .A3(new_n690), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT103), .B(G472), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n643), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n286), .B1(new_n282), .B2(new_n322), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n192), .B(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n603), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n712), .A2(new_n338), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(new_n565), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(G122), .Z(G24));
  AOI21_X1  g553(.A(G902), .B1(new_n311), .B2(new_n312), .ZN(new_n740));
  INV_X1    g554(.A(new_n730), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n661), .B(new_n734), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n705), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n726), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n370), .ZN(G27));
  AOI211_X1 g560(.A(new_n634), .B(new_n604), .C1(new_n524), .C2(new_n521), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n327), .A2(new_n747), .A3(new_n709), .A4(new_n705), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n748), .B2(KEYINPUT104), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n309), .A2(KEYINPUT105), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n309), .A2(KEYINPUT105), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n326), .A2(new_n305), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n565), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n704), .A2(new_n751), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n747), .A2(new_n760), .ZN(new_n761));
  OAI22_X1  g575(.A1(new_n750), .A2(new_n752), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND4_X1  g577(.A1(new_n327), .A2(new_n747), .A3(new_n709), .A4(new_n671), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n699), .A2(new_n328), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n613), .B2(KEYINPUT107), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n613), .B1(new_n630), .B2(new_n631), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n644), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n661), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n766), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n595), .B2(new_n599), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n569), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n595), .A2(KEYINPUT45), .A3(new_n599), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n601), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n601), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n593), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n603), .A3(new_n686), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT106), .Z(new_n785));
  OR2_X1    g599(.A1(new_n774), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n603), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(KEYINPUT47), .A3(new_n603), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n634), .B1(new_n524), .B2(new_n521), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n327), .A2(new_n709), .A3(new_n704), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT108), .ZN(new_n796));
  XOR2_X1   g610(.A(KEYINPUT109), .B(G140), .Z(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G42));
  NOR2_X1   g612(.A1(G952), .A2(G953), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n742), .A2(new_n704), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n747), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n650), .A2(new_n670), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n438), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n699), .A2(KEYINPUT110), .A3(new_n328), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n327), .A2(new_n805), .A3(new_n663), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT110), .B1(new_n793), .B2(new_n804), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n764), .B(new_n802), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n807), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n679), .A3(new_n805), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT111), .A3(new_n764), .A4(new_n802), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n706), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n680), .A2(new_n681), .A3(new_n714), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n679), .B1(new_n816), .B2(new_n801), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n657), .A2(new_n670), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n661), .B(new_n818), .C1(new_n677), .C2(new_n696), .ZN(new_n819));
  INV_X1    g633(.A(new_n729), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n684), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n716), .B1(new_n640), .B2(new_n652), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n726), .A2(new_n725), .B1(new_n729), .B2(new_n737), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n632), .A2(new_n440), .A3(new_n441), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n613), .A2(new_n650), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(new_n826), .A3(new_n612), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n524), .A2(new_n328), .A3(new_n521), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n605), .A4(new_n644), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n606), .A2(new_n664), .A3(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n823), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n814), .A2(new_n762), .A3(new_n822), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n819), .A2(new_n820), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n684), .A2(new_n817), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n800), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n762), .A2(new_n831), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n668), .A2(new_n706), .B1(new_n726), .B2(new_n744), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n673), .B2(new_n683), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n839), .A2(new_n821), .B1(new_n810), .B2(new_n813), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n837), .A2(new_n840), .A3(new_n841), .A4(KEYINPUT53), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n836), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n832), .B2(new_n835), .ZN(new_n846));
  INV_X1    g660(.A(new_n800), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n837), .A2(new_n840), .A3(new_n841), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n843), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT113), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n848), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n836), .A2(new_n842), .A3(new_n843), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n766), .A2(new_n333), .A3(new_n714), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n857), .A2(new_n709), .A3(new_n697), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n613), .A2(new_n632), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n857), .A2(new_n769), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n743), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n858), .A2(new_n859), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(KEYINPUT51), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n790), .B(new_n791), .C1(new_n603), .C2(new_n712), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n731), .A2(new_n734), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n769), .A2(new_n872), .A3(new_n334), .A4(new_n565), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n766), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n700), .A2(new_n634), .A3(new_n715), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n873), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(KEYINPUT50), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n878), .A2(KEYINPUT116), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n877), .A2(KEYINPUT114), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(KEYINPUT116), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n879), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n867), .A2(new_n875), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n868), .A2(new_n874), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n866), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT51), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n861), .A2(new_n565), .A3(new_n758), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT48), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n858), .A2(new_n633), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n893), .B(new_n330), .C1(new_n726), .C2(new_n873), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n887), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n799), .B1(new_n856), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n712), .B(KEYINPUT49), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n565), .A2(new_n328), .A3(new_n603), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n768), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n700), .A2(new_n697), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT119), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n889), .A2(new_n885), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n886), .B(new_n895), .C1(new_n906), .C2(KEYINPUT51), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n850), .B2(new_n855), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n905), .B(new_n902), .C1(new_n908), .C2(new_n799), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n904), .A2(new_n909), .ZN(G75));
  NOR2_X1   g724(.A1(new_n335), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n188), .B1(new_n836), .B2(new_n842), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT56), .B1(new_n913), .B2(G210), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n510), .B(KEYINPUT120), .Z(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT55), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n513), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n912), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n913), .B(KEYINPUT121), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n520), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(G51));
  INV_X1    g737(.A(new_n778), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n836), .A2(new_n842), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n854), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n601), .B(KEYINPUT57), .Z(new_n928));
  AOI21_X1  g742(.A(new_n710), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n924), .A2(new_n919), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n911), .B1(new_n931), .B2(new_n932), .ZN(G54));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n919), .A2(new_n433), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n433), .B1(new_n919), .B2(new_n934), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n911), .ZN(G60));
  NAND2_X1  g751(.A1(new_n624), .A2(new_n626), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  AOI211_X1 g754(.A(new_n938), .B(new_n940), .C1(new_n926), .C2(new_n854), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n850), .A2(new_n855), .A3(new_n942), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n911), .B(new_n941), .C1(new_n938), .C2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n836), .B2(new_n842), .ZN(new_n947));
  INV_X1    g761(.A(new_n660), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n553), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n949), .B(new_n912), .C1(new_n950), .C2(new_n947), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(KEYINPUT123), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(KEYINPUT123), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT124), .Z(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G66));
  INV_X1    g770(.A(new_n337), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n335), .B1(new_n957), .B2(G224), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n824), .A2(new_n830), .ZN(new_n959));
  INV_X1    g773(.A(new_n823), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n961), .B2(new_n335), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n915), .B1(G898), .B2(new_n335), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT125), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  AND2_X1   g779(.A1(new_n839), .A2(new_n702), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n825), .A2(new_n826), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n766), .A2(new_n687), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n709), .A3(new_n327), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n796), .A2(new_n786), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(KEYINPUT62), .B2(new_n967), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n969), .A2(new_n335), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n419), .B(KEYINPUT126), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n275), .B(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n758), .A2(new_n565), .A3(new_n820), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n785), .B1(new_n774), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n838), .B(new_n981), .C1(new_n673), .C2(new_n683), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n762), .A3(new_n796), .A4(new_n764), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n335), .ZN(new_n984));
  INV_X1    g798(.A(new_n978), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n584), .A2(G900), .A3(G953), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n979), .A2(new_n987), .ZN(G72));
  NAND3_X1  g802(.A1(new_n969), .A2(new_n974), .A3(new_n831), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  AOI211_X1 g805(.A(new_n281), .B(new_n276), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n983), .A2(new_n961), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n316), .B1(new_n993), .B2(new_n991), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n316), .A2(new_n991), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n693), .B(new_n995), .C1(new_n846), .C2(new_n848), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n992), .A2(new_n994), .A3(new_n911), .A4(new_n996), .ZN(G57));
endmodule


