//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT94), .ZN(new_n206));
  AOI21_X1  g005(.A(G8gat), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n208), .B2(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n207), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT95), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT91), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT91), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n218), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI211_X1 g022(.A(G29gat), .B(G36gat), .C1(new_n219), .C2(KEYINPUT14), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(new_n222), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT15), .B(new_n216), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(KEYINPUT93), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT92), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n230), .B2(KEYINPUT15), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n231), .C1(KEYINPUT15), .C2(new_n230), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n214), .A2(new_n215), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n215), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n227), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n234), .A2(new_n235), .A3(new_n213), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n203), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(KEYINPUT17), .A3(new_n227), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n211), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n235), .B1(new_n234), .B2(new_n213), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT18), .A4(new_n202), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT11), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n237), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n242), .A3(new_n202), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT96), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n255), .A3(new_n252), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(new_n237), .A3(new_n243), .ZN(new_n258));
  INV_X1    g057(.A(new_n249), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G197gat), .ZN(new_n267));
  INV_X1    g066(.A(G204gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270));
  OAI22_X1  g069(.A1(KEYINPUT22), .A2(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT74), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n273));
  OAI221_X1 g072(.A(new_n273), .B1(new_n266), .B2(KEYINPUT22), .C1(new_n270), .C2(new_n269), .ZN(new_n274));
  XOR2_X1   g073(.A(G211gat), .B(G218gat), .Z(new_n275));
  AND3_X1   g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n272), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n263), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G148gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G141gat), .ZN(new_n282));
  INV_X1    g081(.A(G141gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G148gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n282), .A2(new_n284), .B1(KEYINPUT2), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT78), .A2(G155gat), .A3(G162gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT79), .B1(new_n283), .B2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n281), .A3(G141gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(new_n284), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n285), .B1(new_n289), .B2(KEYINPUT2), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT80), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT80), .B1(new_n297), .B2(new_n298), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n276), .A2(new_n277), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n297), .A2(new_n298), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n292), .B1(new_n307), .B2(new_n299), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n279), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n304), .B1(new_n310), .B2(KEYINPUT29), .ZN(new_n311));
  INV_X1    g110(.A(G228gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n303), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(new_n303), .B2(new_n311), .ZN(new_n316));
  OAI21_X1  g115(.A(G22gat), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n276), .A2(new_n277), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(new_n263), .B2(new_n309), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n308), .B1(new_n278), .B2(new_n279), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n319), .A2(new_n320), .B1(new_n312), .B2(new_n313), .ZN(new_n321));
  INV_X1    g120(.A(G22gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n311), .A3(new_n314), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G78gat), .B(G106gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT31), .ZN(new_n327));
  INV_X1    g126(.A(G50gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT86), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n321), .A2(new_n323), .A3(new_n334), .A4(new_n322), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n324), .A2(KEYINPUT86), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n329), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n330), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G57gat), .B(G85gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(G113gat), .A2(G120gat), .ZN(new_n347));
  INV_X1    g146(.A(G113gat), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n347), .ZN(new_n353));
  AND2_X1   g152(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n355));
  INV_X1    g154(.A(G127gat), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G134gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT66), .B1(new_n358), .B2(G127gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n356), .A3(G134gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n352), .B(new_n353), .C1(new_n357), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n358), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(G127gat), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(new_n359), .A3(new_n361), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n352), .B1(new_n369), .B2(new_n353), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n351), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT68), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n353), .B1(new_n357), .B2(new_n362), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n363), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT68), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n351), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n372), .A2(new_n373), .A3(new_n378), .A4(new_n308), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n371), .A2(new_n302), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n309), .A3(new_n371), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n345), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n307), .A2(new_n299), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n376), .A2(new_n351), .B1(new_n389), .B2(new_n293), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n380), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n302), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n308), .A2(new_n376), .A3(new_n351), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT81), .B1(new_n396), .B2(new_n384), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n378), .A4(new_n308), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n373), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n385), .A3(new_n383), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n399), .B1(new_n398), .B2(new_n402), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n387), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n345), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n392), .B1(new_n391), .B2(KEYINPUT5), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n396), .A2(KEYINPUT81), .A3(new_n384), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n402), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n381), .A2(new_n386), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT84), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n404), .B2(new_n405), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n345), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT6), .B1(new_n414), .B2(new_n387), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(KEYINPUT6), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G190gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(G183gat), .ZN(new_n426));
  INV_X1    g225(.A(G183gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(G190gat), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT24), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(KEYINPUT24), .ZN(new_n430));
  NOR2_X1   g229(.A1(G169gat), .A2(G176gat), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n430), .A2(G190gat), .B1(new_n431), .B2(KEYINPUT23), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n431), .A2(KEYINPUT23), .ZN(new_n433));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n429), .A2(new_n432), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT25), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n433), .A2(new_n434), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(new_n429), .A3(new_n432), .A4(KEYINPUT25), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n431), .A2(KEYINPUT26), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n431), .A2(KEYINPUT26), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n427), .B2(KEYINPUT64), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT64), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(KEYINPUT27), .A3(G183gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n425), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n426), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT28), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(KEYINPUT27), .B(G183gat), .Z(new_n451));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n451), .A2(new_n452), .A3(G190gat), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n441), .B(new_n443), .C1(new_n450), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n440), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n263), .ZN(new_n456));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT75), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n457), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n462), .A2(new_n463), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n304), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(new_n457), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n455), .A2(new_n458), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n318), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G8gat), .B(G36gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G64gat), .ZN(new_n472));
  INV_X1    g271(.A(G92gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n467), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n470), .ZN(new_n479));
  INV_X1    g278(.A(new_n474), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n477), .B1(new_n475), .B2(new_n476), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n340), .B1(new_n424), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n372), .A2(new_n378), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n455), .ZN(new_n488));
  INV_X1    g287(.A(new_n455), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n372), .A3(new_n378), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT33), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G43gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT69), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(G71gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(G71gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G99gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(G99gat), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n502), .ZN(new_n505));
  AOI21_X1  g304(.A(G99gat), .B1(new_n497), .B2(new_n498), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT70), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n508), .A3(new_n502), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(KEYINPUT33), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n510), .A2(KEYINPUT32), .ZN(new_n511));
  INV_X1    g310(.A(new_n491), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n494), .A2(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n488), .A2(new_n486), .A3(new_n490), .ZN(new_n514));
  INV_X1    g313(.A(new_n486), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT34), .B1(new_n515), .B2(KEYINPUT71), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n488), .A2(new_n490), .A3(new_n486), .A4(new_n516), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT73), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n513), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n511), .A2(new_n512), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n504), .B1(new_n491), .B2(new_n493), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n520), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n522), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT72), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n520), .B1(new_n513), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT72), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT36), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT87), .B1(new_n485), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT87), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n482), .A2(new_n483), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n413), .A2(new_n403), .B1(new_n381), .B2(new_n386), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n406), .B(new_n407), .C1(new_n542), .C2(new_n409), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n543), .A2(KEYINPUT84), .B1(KEYINPUT6), .B2(new_n416), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n541), .B1(new_n544), .B2(new_n422), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n539), .B(new_n540), .C1(new_n545), .C2(new_n340), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n543), .A2(KEYINPUT88), .B1(KEYINPUT6), .B2(new_n416), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n419), .A2(new_n420), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550));
  INV_X1    g349(.A(new_n466), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n460), .A2(new_n464), .A3(new_n318), .A4(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n552), .A2(KEYINPUT89), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n318), .B1(new_n468), .B2(new_n469), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n552), .B2(KEYINPUT89), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n550), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n467), .A2(new_n550), .A3(new_n470), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT38), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n480), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n475), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n557), .A2(new_n480), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n479), .A2(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n549), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n340), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n484), .A2(new_n416), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n385), .B1(new_n381), .B2(new_n383), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT39), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n345), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n394), .A2(new_n395), .A3(new_n385), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT39), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT40), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n566), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n538), .A2(new_n546), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n547), .A2(new_n549), .ZN(new_n578));
  INV_X1    g377(.A(new_n530), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n579), .A2(new_n541), .A3(new_n566), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n566), .B1(new_n535), .B2(new_n534), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n424), .A2(new_n583), .A3(new_n484), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n262), .B1(new_n577), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G57gat), .B(G64gat), .Z(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  INV_X1    g388(.A(G71gat), .ZN(new_n590));
  INV_X1    g389(.A(G78gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G71gat), .B(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n594), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n214), .B(new_n215), .C1(new_n599), .C2(new_n598), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G183gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n606), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n264), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n615), .B(new_n473), .C1(new_n616), .C2(KEYINPUT7), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n616), .B2(KEYINPUT7), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT99), .B(new_n619), .C1(new_n615), .C2(new_n473), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n621), .B1(new_n615), .B2(new_n473), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G99gat), .B(G106gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n618), .A2(new_n624), .A3(new_n620), .A4(new_n622), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(KEYINPUT100), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n623), .A2(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(new_n627), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n239), .A2(new_n240), .A3(new_n628), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT101), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n628), .ZN(new_n637));
  AND2_X1   g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n637), .A2(new_n235), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n633), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n642));
  XNOR2_X1  g441(.A(G134gat), .B(G162gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n636), .B1(new_n633), .B2(new_n639), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n641), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n598), .B1(new_n627), .B2(KEYINPUT102), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n630), .B2(new_n631), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n626), .B(new_n627), .C1(KEYINPUT102), .C2(new_n598), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n598), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT10), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n632), .B2(new_n628), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n651), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  INV_X1    g459(.A(new_n651), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G204gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(G176gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n614), .A2(new_n650), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n587), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n424), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n541), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G8gat), .B1(new_n674), .B2(new_n484), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT104), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n682), .A2(new_n687), .A3(new_n683), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n674), .B2(new_n540), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n579), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n674), .B2(new_n691), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n340), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n577), .A2(new_n586), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n650), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n670), .B(KEYINPUT105), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n614), .A2(new_n262), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n530), .A2(new_n484), .A3(new_n340), .A4(new_n581), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n547), .B2(new_n549), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n424), .A2(new_n583), .A3(new_n484), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(KEYINPUT35), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n424), .A2(new_n484), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n537), .B1(new_n708), .B2(new_n566), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n706), .A2(new_n707), .B1(new_n709), .B2(new_n576), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n586), .A2(KEYINPUT106), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n650), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n700), .B(new_n702), .C1(new_n712), .C2(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n696), .B1(new_n713), .B2(new_n424), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n707), .B(new_n582), .C1(new_n584), .C2(new_n585), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n708), .A2(new_n566), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n576), .A3(new_n540), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n706), .A2(new_n707), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n649), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n720), .A2(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n721), .A2(KEYINPUT107), .A3(new_n676), .A4(new_n702), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n714), .A2(G29gat), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n614), .A2(new_n650), .A3(new_n670), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n587), .A2(new_n221), .A3(new_n676), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n723), .A2(new_n729), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1328gat));
  NAND4_X1  g530(.A1(new_n587), .A2(new_n222), .A3(new_n541), .A4(new_n724), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT46), .Z(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n713), .B2(new_n484), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G36gat), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n713), .A2(new_n734), .A3(new_n484), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(G1329gat));
  OAI21_X1  g537(.A(G43gat), .B1(new_n713), .B2(new_n540), .ZN(new_n739));
  INV_X1    g538(.A(G43gat), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n587), .A2(new_n740), .A3(new_n530), .A4(new_n724), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT47), .B1(new_n741), .B2(KEYINPUT110), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1330gat));
  OAI21_X1  g543(.A(G50gat), .B1(new_n713), .B2(new_n340), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n587), .A2(new_n328), .A3(new_n566), .A4(new_n724), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g547(.A1(new_n718), .A2(new_n719), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n614), .A2(new_n262), .A3(new_n650), .A4(new_n701), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n676), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g552(.A1(new_n749), .A2(new_n750), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n484), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  OAI21_X1  g558(.A(KEYINPUT111), .B1(new_n754), .B2(new_n579), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n751), .A2(new_n761), .A3(new_n530), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n590), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n751), .A2(G71gat), .A3(new_n537), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n566), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g567(.A1(new_n612), .A2(new_n613), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n262), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT112), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n649), .B(new_n771), .C1(new_n718), .C2(new_n719), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n710), .A2(new_n711), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n649), .A4(new_n771), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n777), .A2(new_n615), .A3(new_n676), .A4(new_n670), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n771), .A2(new_n670), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n700), .B(new_n779), .C1(new_n712), .C2(KEYINPUT44), .ZN(new_n780));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780), .B2(new_n424), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n774), .A2(new_n783), .A3(new_n776), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n772), .A2(KEYINPUT113), .A3(new_n773), .ZN(new_n785));
  INV_X1    g584(.A(new_n701), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n786), .A2(G92gat), .A3(new_n484), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n780), .B2(new_n484), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n772), .A2(new_n773), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n712), .B2(new_n771), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n796));
  NAND3_X1  g595(.A1(new_n789), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n791), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n788), .B2(new_n789), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n789), .A2(new_n795), .A3(new_n796), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(G1337gat));
  NAND4_X1  g602(.A1(new_n777), .A2(new_n500), .A3(new_n530), .A4(new_n670), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n780), .A2(new_n540), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n500), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT116), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n721), .A2(new_n566), .A3(new_n779), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n786), .A2(G106gat), .A3(new_n340), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n784), .A2(new_n785), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n777), .A2(new_n810), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g614(.A(new_n657), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n637), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n661), .C1(KEYINPUT10), .C2(new_n660), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(KEYINPUT54), .A3(new_n659), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n651), .C1(new_n655), .C2(new_n658), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n667), .A4(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n668), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n819), .A2(new_n667), .A3(new_n821), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n823), .B1(new_n822), .B2(new_n668), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT118), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n822), .A2(new_n668), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n833), .A3(new_n827), .A4(new_n824), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n261), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n233), .A2(new_n236), .A3(new_n203), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n202), .B1(new_n241), .B2(new_n242), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n248), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n257), .A2(new_n670), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n649), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n649), .A2(new_n257), .A3(new_n838), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n830), .A2(new_n841), .A3(new_n834), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n769), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n672), .A2(new_n261), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n424), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n580), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n348), .A3(new_n262), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n583), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n261), .A3(new_n484), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n852), .B2(new_n348), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n484), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n349), .B1(new_n854), .B2(new_n671), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n701), .A2(G120gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT119), .ZN(G1341gat));
  OAI21_X1  g657(.A(G127gat), .B1(new_n848), .B2(new_n769), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n614), .A2(new_n356), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n854), .B2(new_n860), .ZN(G1342gat));
  NAND2_X1  g660(.A1(new_n484), .A2(new_n649), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n851), .A2(new_n366), .A3(new_n367), .A4(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n848), .B2(new_n650), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NOR3_X1   g668(.A1(new_n424), .A2(new_n537), .A3(new_n541), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT121), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n566), .A2(KEYINPUT57), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n825), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n831), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n261), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(new_n839), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n877), .B2(new_n839), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n650), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n614), .B1(new_n881), .B2(new_n842), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n873), .B1(new_n882), .B2(new_n845), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT125), .B(new_n873), .C1(new_n882), .C2(new_n845), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n844), .A2(new_n846), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n566), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n885), .B(new_n886), .C1(new_n888), .C2(KEYINPUT122), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n261), .B(new_n871), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G141gat), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n847), .A2(new_n566), .A3(new_n540), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(new_n283), .A3(new_n261), .A4(new_n484), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n892), .B(new_n894), .C1(new_n897), .C2(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1344gat));
  OR2_X1    g700(.A1(new_n889), .A2(new_n890), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n871), .A2(new_n670), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n893), .A2(new_n484), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT59), .B1(new_n906), .B2(new_n671), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n281), .ZN(new_n908));
  INV_X1    g707(.A(new_n881), .ZN(new_n909));
  INV_X1    g708(.A(new_n841), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(new_n829), .A3(new_n828), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n769), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n846), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n566), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n872), .B1(new_n844), .B2(new_n846), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT59), .B(G148gat), .C1(new_n916), .C2(new_n903), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n905), .A2(new_n908), .A3(new_n917), .ZN(G1345gat));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n871), .ZN(new_n919));
  OAI21_X1  g718(.A(G155gat), .B1(new_n919), .B2(new_n769), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n769), .A2(G155gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n906), .B2(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n919), .B2(new_n650), .ZN(new_n923));
  INV_X1    g722(.A(G162gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n893), .A2(new_n924), .A3(new_n864), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1347gat));
  AOI21_X1  g725(.A(new_n676), .B1(new_n844), .B2(new_n846), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(new_n541), .A3(new_n340), .A4(new_n530), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n246), .A3(new_n262), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n583), .A2(new_n541), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n261), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n929), .A2(new_n933), .ZN(G1348gat));
  INV_X1    g733(.A(new_n932), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n935), .A2(G176gat), .A3(new_n671), .ZN(new_n936));
  OAI21_X1  g735(.A(G176gat), .B1(new_n928), .B2(new_n786), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n928), .B2(new_n769), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n769), .A2(new_n451), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n941), .B(new_n942), .Z(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n928), .B2(new_n650), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n425), .A3(new_n649), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  AND4_X1   g746(.A1(new_n541), .A2(new_n927), .A3(new_n566), .A4(new_n540), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n261), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n540), .A2(new_n541), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(new_n676), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n916), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n262), .A2(new_n267), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n268), .A3(new_n670), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT62), .Z(new_n957));
  NOR3_X1   g756(.A1(new_n916), .A2(new_n786), .A3(new_n952), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n268), .B2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n264), .A3(new_n614), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n953), .A2(new_n614), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  AOI21_X1  g763(.A(G218gat), .B1(new_n948), .B2(new_n649), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n650), .A2(new_n265), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n953), .B2(new_n966), .ZN(G1355gat));
endmodule


