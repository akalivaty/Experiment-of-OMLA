

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n315), .B(n314), .ZN(n537) );
  XNOR2_X1 U326 ( .A(n378), .B(n319), .ZN(n323) );
  XNOR2_X1 U327 ( .A(n371), .B(n370), .ZN(n486) );
  XNOR2_X1 U328 ( .A(n449), .B(n369), .ZN(n370) );
  XNOR2_X1 U329 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n465) );
  XNOR2_X1 U330 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U331 ( .A1(n540), .A2(n397), .ZN(n398) );
  XNOR2_X1 U332 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U333 ( .A(n380), .B(n379), .ZN(n381) );
  INV_X1 U334 ( .A(G204GAT), .ZN(n379) );
  NOR2_X1 U335 ( .A1(n537), .A2(n489), .ZN(n574) );
  XNOR2_X1 U336 ( .A(n335), .B(n334), .ZN(n573) );
  XOR2_X1 U337 ( .A(n438), .B(n376), .Z(n293) );
  XOR2_X1 U338 ( .A(G78GAT), .B(n404), .Z(n294) );
  AND2_X1 U339 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U340 ( .A(KEYINPUT112), .B(n458), .Z(n296) );
  NOR2_X1 U341 ( .A1(n487), .A2(n555), .ZN(n587) );
  INV_X1 U342 ( .A(KEYINPUT25), .ZN(n389) );
  XNOR2_X1 U343 ( .A(n389), .B(KEYINPUT95), .ZN(n390) );
  INV_X1 U344 ( .A(KEYINPUT71), .ZN(n443) );
  INV_X1 U345 ( .A(G106GAT), .ZN(n317) );
  XNOR2_X1 U346 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U347 ( .A(n402), .B(n295), .ZN(n360) );
  XNOR2_X1 U348 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U349 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U350 ( .A(n446), .B(n445), .ZN(n447) );
  NOR2_X1 U351 ( .A1(n537), .A2(n554), .ZN(n538) );
  XNOR2_X1 U352 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U353 ( .A1(n475), .A2(n417), .ZN(n418) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n315) );
  INV_X1 U356 ( .A(G218GAT), .ZN(n476) );
  XNOR2_X1 U357 ( .A(KEYINPUT114), .B(n541), .ZN(n550) );
  INV_X1 U358 ( .A(G43GAT), .ZN(n482) );
  XNOR2_X1 U359 ( .A(KEYINPUT38), .B(n481), .ZN(n513) );
  XNOR2_X1 U360 ( .A(n476), .B(KEYINPUT62), .ZN(n477) );
  XNOR2_X1 U361 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U362 ( .A(n317), .B(KEYINPUT44), .ZN(n454) );
  XNOR2_X1 U363 ( .A(n451), .B(KEYINPUT108), .ZN(n452) );
  XNOR2_X1 U364 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U365 ( .A(n478), .B(n477), .ZN(G1355GAT) );
  XNOR2_X1 U366 ( .A(n493), .B(n492), .ZN(G1349GAT) );
  XNOR2_X1 U367 ( .A(n453), .B(n452), .ZN(G1338GAT) );
  XOR2_X1 U368 ( .A(G127GAT), .B(G134GAT), .Z(n298) );
  XNOR2_X1 U369 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n297) );
  XNOR2_X1 U370 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U371 ( .A(G113GAT), .B(n299), .Z(n344) );
  XNOR2_X1 U372 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n300) );
  XNOR2_X1 U373 ( .A(n300), .B(KEYINPUT17), .ZN(n301) );
  XOR2_X1 U374 ( .A(n301), .B(KEYINPUT81), .Z(n303) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U376 ( .A(n303), .B(n302), .ZN(n386) );
  XNOR2_X1 U377 ( .A(n344), .B(n386), .ZN(n313) );
  XOR2_X1 U378 ( .A(G71GAT), .B(G183GAT), .Z(n305) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G176GAT), .ZN(n304) );
  XNOR2_X1 U380 ( .A(n305), .B(n304), .ZN(n307) );
  XOR2_X1 U381 ( .A(G43GAT), .B(G190GAT), .Z(n306) );
  XNOR2_X1 U382 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U383 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n309) );
  XNOR2_X1 U384 ( .A(G15GAT), .B(KEYINPUT79), .ZN(n308) );
  XNOR2_X1 U385 ( .A(n309), .B(n308), .ZN(n310) );
  NAND2_X1 U386 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U388 ( .A(n316), .B(KEYINPUT77), .ZN(n378) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XOR2_X1 U390 ( .A(KEYINPUT76), .B(KEYINPUT65), .Z(n321) );
  XNOR2_X1 U391 ( .A(KEYINPUT75), .B(KEYINPUT9), .ZN(n320) );
  XNOR2_X1 U392 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U393 ( .A(n323), .B(n322), .Z(n329) );
  XOR2_X1 U394 ( .A(G29GAT), .B(G43GAT), .Z(n325) );
  XNOR2_X1 U395 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n324) );
  XNOR2_X1 U396 ( .A(n325), .B(n324), .ZN(n428) );
  XOR2_X1 U397 ( .A(KEYINPUT73), .B(G92GAT), .Z(n327) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G85GAT), .ZN(n326) );
  XNOR2_X1 U399 ( .A(n327), .B(n326), .ZN(n442) );
  XNOR2_X1 U400 ( .A(n428), .B(n442), .ZN(n328) );
  XNOR2_X1 U401 ( .A(n329), .B(n328), .ZN(n335) );
  XNOR2_X1 U402 ( .A(G50GAT), .B(G162GAT), .ZN(n330) );
  XNOR2_X1 U403 ( .A(n330), .B(KEYINPUT74), .ZN(n368) );
  XOR2_X1 U404 ( .A(KEYINPUT10), .B(n368), .Z(n332) );
  XNOR2_X1 U405 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n331) );
  XNOR2_X1 U406 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U407 ( .A(G134GAT), .B(n333), .ZN(n334) );
  XOR2_X1 U408 ( .A(KEYINPUT36), .B(n573), .Z(n475) );
  XOR2_X1 U409 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n337) );
  XNOR2_X1 U410 ( .A(G141GAT), .B(KEYINPUT84), .ZN(n336) );
  XNOR2_X1 U411 ( .A(n337), .B(n336), .ZN(n357) );
  XOR2_X1 U412 ( .A(G85GAT), .B(n357), .Z(n339) );
  NAND2_X1 U413 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U414 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U415 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n341) );
  XNOR2_X1 U416 ( .A(KEYINPUT87), .B(KEYINPUT1), .ZN(n340) );
  XNOR2_X1 U417 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U418 ( .A(n343), .B(n342), .Z(n346) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(n344), .ZN(n345) );
  XNOR2_X1 U420 ( .A(n346), .B(n345), .ZN(n354) );
  XOR2_X1 U421 ( .A(G148GAT), .B(G57GAT), .Z(n348) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(G155GAT), .ZN(n347) );
  XNOR2_X1 U423 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U424 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n350) );
  XNOR2_X1 U425 ( .A(G162GAT), .B(KEYINPUT4), .ZN(n349) );
  XNOR2_X1 U426 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U427 ( .A(n352), .B(n351), .Z(n353) );
  XNOR2_X1 U428 ( .A(n354), .B(n353), .ZN(n534) );
  XOR2_X1 U429 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n356) );
  XNOR2_X1 U430 ( .A(G197GAT), .B(G218GAT), .ZN(n355) );
  XNOR2_X1 U431 ( .A(n356), .B(n355), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n357), .B(n373), .ZN(n363) );
  XOR2_X1 U433 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n359) );
  XNOR2_X1 U434 ( .A(G211GAT), .B(KEYINPUT23), .ZN(n358) );
  XNOR2_X1 U435 ( .A(n359), .B(n358), .ZN(n361) );
  XOR2_X1 U436 ( .A(G22GAT), .B(G155GAT), .Z(n402) );
  XNOR2_X1 U437 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U438 ( .A(n364), .B(KEYINPUT85), .Z(n371) );
  XOR2_X1 U439 ( .A(KEYINPUT72), .B(G78GAT), .Z(n366) );
  XNOR2_X1 U440 ( .A(G148GAT), .B(G106GAT), .ZN(n365) );
  XNOR2_X1 U441 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U442 ( .A(G204GAT), .B(n367), .Z(n449) );
  XNOR2_X1 U443 ( .A(n368), .B(KEYINPUT24), .ZN(n369) );
  XNOR2_X1 U444 ( .A(G8GAT), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U445 ( .A(n372), .B(G211GAT), .ZN(n404) );
  XNOR2_X1 U446 ( .A(n373), .B(n404), .ZN(n384) );
  XOR2_X1 U447 ( .A(G176GAT), .B(G64GAT), .Z(n438) );
  XOR2_X1 U448 ( .A(KEYINPUT93), .B(KEYINPUT90), .Z(n375) );
  XNOR2_X1 U449 ( .A(G92GAT), .B(KEYINPUT91), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n375), .B(n374), .ZN(n376) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U452 ( .A(n293), .B(n377), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n378), .B(KEYINPUT92), .ZN(n380) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n470) );
  NOR2_X1 U456 ( .A1(n537), .A2(n470), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n387), .B(KEYINPUT94), .ZN(n388) );
  NOR2_X1 U458 ( .A1(n486), .A2(n388), .ZN(n391) );
  NAND2_X1 U459 ( .A1(n534), .A2(n392), .ZN(n395) );
  XNOR2_X1 U460 ( .A(KEYINPUT27), .B(n470), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n486), .A2(n537), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n393), .B(KEYINPUT26), .ZN(n555) );
  NOR2_X1 U463 ( .A1(n396), .A2(n555), .ZN(n394) );
  NOR2_X1 U464 ( .A1(n395), .A2(n394), .ZN(n400) );
  XOR2_X1 U465 ( .A(KEYINPUT28), .B(n486), .Z(n525) );
  INV_X1 U466 ( .A(n525), .ZN(n540) );
  INV_X1 U467 ( .A(n396), .ZN(n535) );
  NAND2_X1 U468 ( .A1(n537), .A2(n535), .ZN(n397) );
  NOR2_X1 U469 ( .A1(n398), .A2(n534), .ZN(n399) );
  NOR2_X1 U470 ( .A1(n400), .A2(n399), .ZN(n401) );
  XOR2_X1 U471 ( .A(KEYINPUT96), .B(n401), .Z(n497) );
  XNOR2_X1 U472 ( .A(G127GAT), .B(G64GAT), .ZN(n403) );
  XOR2_X1 U473 ( .A(n403), .B(n402), .Z(n415) );
  NAND2_X1 U474 ( .A1(G231GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n294), .B(n405), .ZN(n409) );
  XOR2_X1 U476 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n407) );
  XNOR2_X1 U477 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U479 ( .A(n409), .B(n408), .Z(n413) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n410), .B(G15GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(G71GAT), .B(G57GAT), .ZN(n411) );
  XNOR2_X1 U483 ( .A(n411), .B(KEYINPUT13), .ZN(n439) );
  XNOR2_X1 U484 ( .A(n426), .B(n439), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X2 U486 ( .A(n415), .B(n414), .Z(n586) );
  NOR2_X1 U487 ( .A1(n497), .A2(n586), .ZN(n416) );
  XOR2_X1 U488 ( .A(KEYINPUT100), .B(n416), .Z(n417) );
  XOR2_X1 U489 ( .A(KEYINPUT37), .B(n418), .Z(n480) );
  XOR2_X1 U490 ( .A(G22GAT), .B(G8GAT), .Z(n420) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U493 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n422) );
  XNOR2_X1 U494 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n421) );
  XNOR2_X1 U495 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U496 ( .A(n424), .B(n423), .ZN(n435) );
  XNOR2_X1 U497 ( .A(G113GAT), .B(G36GAT), .ZN(n425) );
  XNOR2_X1 U498 ( .A(n425), .B(G50GAT), .ZN(n427) );
  XOR2_X1 U499 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U500 ( .A(n428), .B(KEYINPUT67), .Z(n430) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U502 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U503 ( .A(n431), .B(G141GAT), .ZN(n432) );
  XNOR2_X1 U504 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U505 ( .A(n435), .B(n434), .Z(n479) );
  INV_X1 U506 ( .A(n479), .ZN(n579) );
  XOR2_X1 U507 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n437) );
  XNOR2_X1 U508 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n436) );
  XNOR2_X1 U509 ( .A(n437), .B(n436), .ZN(n448) );
  XOR2_X1 U510 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U512 ( .A(n441), .B(n440), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n442), .B(KEYINPUT33), .ZN(n444) );
  XNOR2_X1 U514 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X2 U515 ( .A(n450), .B(n449), .Z(n582) );
  XNOR2_X1 U516 ( .A(KEYINPUT41), .B(n582), .ZN(n459) );
  NOR2_X1 U517 ( .A1(n579), .A2(n459), .ZN(n517) );
  NAND2_X1 U518 ( .A1(n480), .A2(n517), .ZN(n531) );
  NOR2_X1 U519 ( .A1(n537), .A2(n531), .ZN(n453) );
  INV_X1 U520 ( .A(G99GAT), .ZN(n451) );
  NOR2_X1 U521 ( .A1(n525), .A2(n531), .ZN(n455) );
  XNOR2_X1 U522 ( .A(n455), .B(n454), .ZN(G1339GAT) );
  INV_X1 U523 ( .A(n586), .ZN(n494) );
  NOR2_X1 U524 ( .A1(n494), .A2(n475), .ZN(n456) );
  XOR2_X1 U525 ( .A(KEYINPUT45), .B(n456), .Z(n457) );
  NOR2_X1 U526 ( .A1(n582), .A2(n457), .ZN(n458) );
  OR2_X1 U527 ( .A1(n579), .A2(n296), .ZN(n468) );
  XOR2_X1 U528 ( .A(KEYINPUT109), .B(n586), .Z(n569) );
  NOR2_X1 U529 ( .A1(n459), .A2(n479), .ZN(n460) );
  XNOR2_X1 U530 ( .A(n460), .B(KEYINPUT46), .ZN(n461) );
  NOR2_X1 U531 ( .A1(n569), .A2(n461), .ZN(n462) );
  XNOR2_X1 U532 ( .A(n462), .B(KEYINPUT110), .ZN(n464) );
  INV_X1 U533 ( .A(n573), .ZN(n463) );
  NAND2_X1 U534 ( .A1(n464), .A2(n463), .ZN(n466) );
  AND2_X1 U535 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U536 ( .A(n469), .B(KEYINPUT48), .ZN(n533) );
  NOR2_X1 U537 ( .A1(n470), .A2(n533), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n471), .B(KEYINPUT54), .ZN(n472) );
  NAND2_X1 U539 ( .A1(n472), .A2(n534), .ZN(n473) );
  XNOR2_X1 U540 ( .A(n473), .B(KEYINPUT64), .ZN(n487) );
  INV_X1 U541 ( .A(n587), .ZN(n474) );
  NOR2_X1 U542 ( .A1(n475), .A2(n474), .ZN(n478) );
  NOR2_X1 U543 ( .A1(n479), .A2(n582), .ZN(n498) );
  NAND2_X1 U544 ( .A1(n480), .A2(n498), .ZN(n481) );
  NOR2_X1 U545 ( .A1(n537), .A2(n513), .ZN(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(G1330GAT) );
  NOR2_X1 U548 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT55), .ZN(n489) );
  INV_X1 U550 ( .A(n459), .ZN(n560) );
  NAND2_X1 U551 ( .A1(n574), .A2(n560), .ZN(n493) );
  XOR2_X1 U552 ( .A(G176GAT), .B(KEYINPUT56), .Z(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n490) );
  NOR2_X1 U554 ( .A1(n573), .A2(n494), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(n495), .Z(n496) );
  NOR2_X1 U556 ( .A1(n497), .A2(n496), .ZN(n516) );
  NAND2_X1 U557 ( .A1(n498), .A2(n516), .ZN(n506) );
  NOR2_X1 U558 ( .A1(n534), .A2(n506), .ZN(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NOR2_X1 U562 ( .A1(n470), .A2(n506), .ZN(n502) );
  XOR2_X1 U563 ( .A(G8GAT), .B(n502), .Z(G1325GAT) );
  NOR2_X1 U564 ( .A1(n537), .A2(n506), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G15GAT), .B(n505), .ZN(G1326GAT) );
  NOR2_X1 U568 ( .A1(n525), .A2(n506), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1327GAT) );
  NOR2_X1 U571 ( .A1(n513), .A2(n534), .ZN(n510) );
  XNOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  NOR2_X1 U574 ( .A1(n513), .A2(n470), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1329GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n525), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n516), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n534), .A2(n524), .ZN(n519) );
  XNOR2_X1 U582 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n520), .Z(G1332GAT) );
  NOR2_X1 U585 ( .A1(n470), .A2(n524), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1333GAT) );
  NOR2_X1 U588 ( .A1(n537), .A2(n524), .ZN(n523) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G78GAT), .B(n528), .ZN(G1335GAT) );
  NOR2_X1 U594 ( .A1(n534), .A2(n531), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1336GAT) );
  NOR2_X1 U597 ( .A1(n470), .A2(n531), .ZN(n532) );
  XOR2_X1 U598 ( .A(G92GAT), .B(n532), .Z(G1337GAT) );
  XOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT115), .Z(n543) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n554) );
  XNOR2_X1 U602 ( .A(n538), .B(KEYINPUT113), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n579), .A2(n550), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U607 ( .A1(n550), .A2(n560), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n548) );
  NAND2_X1 U611 ( .A1(n550), .A2(n569), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n552) );
  NAND2_X1 U615 ( .A1(n573), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n579), .A2(n565), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n558) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT119), .B(n559), .Z(n562) );
  NAND2_X1 U625 ( .A1(n565), .A2(n560), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(G155GAT), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n586), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n573), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n574), .A2(n579), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n574), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT124), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT58), .B(n572), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1351GAT) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT60), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(n578), .Z(n581) );
  NAND2_X1 U645 ( .A1(n587), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
endmodule

