//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT74), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n192));
  OAI211_X1 g006(.A(G146), .B(new_n190), .C1(new_n192), .C2(new_n188), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  INV_X1    g012(.A(G110), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n197), .A2(new_n198), .A3(new_n199), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n195), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n202), .A2(new_n205), .B1(new_n206), .B2(new_n191), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n193), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G137), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n209), .B(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n187), .A2(G140), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT16), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n188), .B1(new_n216), .B2(new_n189), .ZN(new_n217));
  INV_X1    g031(.A(new_n190), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n206), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n219), .A2(new_n193), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n197), .A2(new_n201), .A3(new_n198), .ZN(new_n221));
  OAI22_X1  g035(.A1(new_n221), .A2(new_n199), .B1(new_n203), .B2(new_n204), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n208), .B(new_n212), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n212), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n219), .B2(new_n193), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n193), .A2(new_n207), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT73), .B(G217), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(G234), .B2(new_n230), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n228), .A2(G902), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n227), .A3(new_n230), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n223), .A2(new_n227), .A3(KEYINPUT25), .A4(new_n230), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n237), .B2(new_n231), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .A3(G134), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G137), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT65), .B(new_n246), .C1(new_n242), .C2(G137), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(G134), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT65), .B1(new_n249), .B2(new_n246), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n244), .B(new_n245), .C1(new_n248), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n243), .A3(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(G131), .C1(new_n252), .C2(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n206), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT1), .B1(new_n258), .B2(G146), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n258), .C2(G146), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(G128), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(new_n259), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n255), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n244), .B1(new_n248), .B2(new_n250), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G131), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n277), .B2(new_n251), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n200), .A2(G116), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G119), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT2), .B(G113), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT28), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n255), .B2(new_n267), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n272), .A2(new_n274), .ZN(new_n290));
  INV_X1    g104(.A(new_n251), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n246), .B1(new_n242), .B2(G137), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n247), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n245), .B1(new_n295), .B2(new_n244), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n290), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n264), .A2(G128), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT67), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n266), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n260), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(KEYINPUT68), .A3(new_n251), .A4(new_n254), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n289), .A2(new_n297), .A3(new_n303), .A4(new_n286), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n279), .B2(new_n286), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n287), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G237), .ZN(new_n311));
  AOI21_X1  g125(.A(G953), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G210), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT27), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G101), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n289), .A2(new_n297), .A3(new_n303), .A4(KEYINPUT30), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n268), .B2(new_n278), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n320), .A3(new_n285), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n321), .A2(new_n304), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT31), .A4(new_n316), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n316), .A4(new_n304), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n317), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT32), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n325), .A2(new_n326), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n325), .A2(new_n326), .ZN(new_n333));
  OAI22_X1  g147(.A1(new_n332), .A2(new_n333), .B1(new_n316), .B2(new_n307), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT32), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n329), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n307), .A2(new_n316), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n321), .A2(new_n304), .ZN(new_n340));
  INV_X1    g154(.A(new_n316), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n287), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n297), .B1(new_n267), .B2(new_n255), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n285), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT72), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n289), .A2(new_n297), .A3(new_n303), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n285), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n352), .B2(new_n304), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n316), .A2(KEYINPUT29), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n343), .B(new_n230), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G472), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n239), .B1(new_n337), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n309), .A2(new_n311), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT85), .A2(G143), .ZN(new_n360));
  OAI21_X1  g174(.A(G214), .B1(KEYINPUT85), .B2(G143), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n210), .A2(new_n359), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n360), .B1(new_n312), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n245), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT17), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n210), .A3(new_n362), .ZN(new_n367));
  INV_X1    g181(.A(new_n360), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n312), .A2(new_n360), .A3(new_n362), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(G131), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n363), .A2(new_n364), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT17), .A4(G131), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n369), .A2(KEYINPUT17), .A3(G131), .A4(new_n370), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT89), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n372), .A2(new_n375), .A3(new_n220), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n191), .B(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n369), .A2(new_n370), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n381), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT86), .B1(new_n373), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n369), .A2(KEYINPUT86), .A3(new_n383), .A4(new_n370), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n378), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n217), .A2(new_n218), .A3(new_n206), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n214), .A2(new_n215), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT19), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n191), .A2(KEYINPUT19), .ZN(new_n396));
  AOI21_X1  g210(.A(G146), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT87), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n365), .A2(new_n371), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n206), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n193), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n387), .A2(KEYINPUT88), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n390), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT88), .B1(new_n387), .B2(new_n404), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n391), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NOR2_X1   g224(.A1(G475), .A2(G902), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n409), .A2(KEYINPUT90), .A3(new_n410), .A4(new_n411), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n378), .A2(new_n387), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n406), .ZN(new_n420));
  AOI211_X1 g234(.A(KEYINPUT92), .B(new_n390), .C1(new_n378), .C2(new_n387), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n391), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n230), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(KEYINPUT93), .A3(new_n230), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT91), .B(G475), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n258), .A2(G128), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n194), .A2(G143), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G134), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n435), .A3(new_n242), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n281), .A2(KEYINPUT14), .A3(G122), .ZN(new_n440));
  XOR2_X1   g254(.A(G116), .B(G122), .Z(new_n441));
  OAI211_X1 g255(.A(G107), .B(new_n440), .C1(new_n441), .C2(KEYINPUT14), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G122), .ZN(new_n443));
  INV_X1    g257(.A(G107), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n439), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(G107), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT95), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n445), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n448), .B2(new_n438), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT13), .B1(new_n258), .B2(G128), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT94), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n436), .B1(KEYINPUT13), .B2(new_n434), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n242), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n446), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT9), .B(G234), .Z(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT75), .ZN(new_n457));
  INV_X1    g271(.A(new_n229), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n210), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n446), .C1(new_n454), .C2(new_n450), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n432), .B1(new_n463), .B2(new_n230), .ZN(new_n464));
  AOI211_X1 g278(.A(G902), .B(new_n431), .C1(new_n460), .C2(new_n462), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(G234), .A2(G237), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(G952), .A3(new_n210), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(G902), .A3(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n417), .A2(new_n429), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G221), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n457), .B2(new_n230), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n444), .A3(G104), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n389), .A2(G107), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G101), .ZN(new_n483));
  INV_X1    g297(.A(G101), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(new_n480), .A3(new_n484), .A4(new_n481), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n487), .A3(G101), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n290), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n389), .A2(G107), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n444), .A2(G104), .ZN(new_n491));
  OAI21_X1  g305(.A(G101), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n485), .A2(new_n492), .A3(KEYINPUT10), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n302), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n261), .A2(G128), .B1(new_n257), .B2(new_n259), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n485), .B(new_n492), .C1(new_n495), .C2(new_n260), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT10), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n277), .A2(new_n251), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n500), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n302), .A2(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n489), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n210), .A2(G227), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT76), .ZN(new_n507));
  XOR2_X1   g321(.A(G110), .B(G140), .Z(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n485), .A2(new_n492), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n496), .B1(new_n302), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n500), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT12), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n502), .A3(new_n489), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n500), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n509), .B(KEYINPUT77), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n505), .A2(new_n509), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G469), .B1(new_n520), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n509), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n501), .B2(new_n504), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n514), .A2(new_n515), .A3(new_n509), .A4(new_n517), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G469), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n230), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n477), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G210), .B1(G237), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT83), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT82), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n283), .A2(new_n284), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n510), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G113), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n281), .A2(G119), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT5), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT5), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT78), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n539), .A2(KEYINPUT78), .A3(new_n540), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G122), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n486), .A2(new_n285), .A3(new_n488), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n300), .A2(new_n187), .A3(new_n301), .ZN(new_n547));
  INV_X1    g361(.A(new_n269), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n273), .A2(new_n548), .A3(new_n270), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n269), .B1(new_n266), .B2(new_n271), .ZN(new_n550));
  OAI21_X1  g364(.A(G125), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n210), .A2(G224), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n542), .A2(new_n541), .B1(new_n283), .B2(new_n284), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT79), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n540), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n540), .A2(new_n558), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n539), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n557), .A2(new_n510), .B1(new_n535), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n544), .B(KEYINPUT8), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n546), .B(new_n556), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT80), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT7), .B1(new_n554), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n566), .B2(new_n554), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n547), .A2(new_n551), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n547), .A2(new_n551), .A3(KEYINPUT81), .A4(new_n568), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n533), .B(new_n230), .C1(new_n565), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n543), .A2(new_n545), .ZN(new_n575));
  INV_X1    g389(.A(new_n544), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n552), .B(new_n555), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT6), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n561), .A2(new_n535), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n539), .A2(new_n540), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n539), .A2(KEYINPUT78), .A3(new_n540), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n534), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n589), .B2(new_n511), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n563), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n571), .A2(new_n572), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n546), .A4(new_n556), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n533), .B1(new_n593), .B2(new_n230), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n532), .B1(new_n583), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n230), .B1(new_n565), .B2(new_n573), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(new_n531), .A3(new_n582), .A4(new_n574), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G214), .B1(G237), .B2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT84), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(KEYINPUT84), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n358), .A2(new_n475), .A3(new_n528), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  AOI21_X1  g421(.A(G478), .B1(new_n463), .B2(new_n230), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n463), .B1(KEYINPUT96), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(KEYINPUT96), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n610), .B(new_n611), .Z(new_n612));
  NOR2_X1   g426(.A1(new_n430), .A2(G902), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n417), .B2(new_n429), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n334), .B2(new_n230), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n328), .A2(new_n330), .ZN(new_n618));
  NAND2_X1  g432(.A1(G469), .A2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n518), .A2(new_n519), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n499), .A2(new_n500), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n515), .A3(new_n509), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(G469), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n527), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n477), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n238), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n617), .A2(new_n618), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n600), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n597), .A2(new_n582), .A3(new_n574), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(new_n529), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n597), .A2(new_n530), .A3(new_n582), .A4(new_n574), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n473), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n615), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n391), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n193), .A2(new_n401), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n638), .A2(KEYINPUT87), .B1(new_n365), .B2(new_n371), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n369), .A2(new_n383), .A3(new_n370), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT86), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n385), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n639), .A2(new_n403), .B1(new_n643), .B2(new_n382), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n390), .B1(new_n644), .B2(KEYINPUT88), .ZN(new_n645));
  INV_X1    g459(.A(new_n408), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n637), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n411), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT20), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(KEYINPUT97), .A3(new_n412), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(KEYINPUT20), .C1(new_n647), .C2(new_n648), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n650), .A2(new_n466), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n429), .A2(KEYINPUT98), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n427), .B1(new_n423), .B2(new_n424), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n426), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n473), .B(KEYINPUT99), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n653), .A2(new_n654), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n632), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n656), .A2(new_n425), .A3(new_n426), .A4(new_n428), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n656), .B1(new_n655), .B2(new_n426), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(KEYINPUT100), .A3(new_n653), .A4(new_n658), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n662), .B1(new_n661), .B2(new_n666), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n627), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NOR2_X1   g485(.A1(new_n617), .A2(new_n618), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n237), .A2(new_n231), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n225), .A2(new_n226), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n677), .B(new_n230), .C1(G234), .C2(new_n229), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n528), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n475), .A2(new_n605), .A3(new_n672), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NAND4_X1  g497(.A1(new_n528), .A2(new_n630), .A3(new_n631), .A4(new_n679), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n337), .B2(new_n357), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n470), .A2(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n468), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n685), .A2(new_n665), .A3(new_n653), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XNOR2_X1  g503(.A(new_n687), .B(KEYINPUT39), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n528), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT102), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT40), .Z(new_n693));
  NOR2_X1   g507(.A1(new_n340), .A2(new_n341), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n316), .B1(new_n352), .B2(new_n304), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n230), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n337), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n599), .B(KEYINPUT38), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n417), .A2(new_n429), .ZN(new_n700));
  INV_X1    g514(.A(new_n679), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n600), .A3(new_n466), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n693), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  NAND3_X1  g519(.A1(new_n685), .A2(new_n615), .A3(new_n687), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  AOI21_X1  g521(.A(G902), .B1(new_n523), .B2(new_n524), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n526), .A2(KEYINPUT103), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n625), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n358), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n615), .A2(new_n633), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  INV_X1    g532(.A(new_n714), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n667), .B2(new_n668), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND2_X1  g535(.A1(new_n337), .A2(new_n357), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n632), .A2(new_n701), .A3(new_n712), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n475), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND3_X1  g539(.A1(new_n630), .A2(new_n466), .A3(new_n631), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n417), .B2(new_n429), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n324), .A2(new_n327), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n341), .B1(new_n350), .B2(new_n353), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n330), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n617), .A2(new_n730), .A3(new_n239), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n727), .A2(new_n731), .A3(new_n658), .A4(new_n713), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR3_X1   g547(.A1(new_n617), .A2(new_n730), .A3(new_n701), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n632), .A2(new_n712), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n615), .A2(new_n734), .A3(new_n687), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n619), .B(KEYINPUT104), .Z(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n708), .B2(new_n526), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n622), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n621), .A2(new_n515), .A3(KEYINPUT105), .A4(new_n509), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(G469), .A3(new_n620), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT106), .B1(new_n747), .B2(new_n625), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n749), .B(new_n477), .C1(new_n741), .C2(new_n746), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n595), .A2(new_n600), .A3(new_n598), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n615), .A3(new_n687), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n722), .A2(new_n238), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n738), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n687), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n756), .B(new_n614), .C1(new_n417), .C2(new_n429), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n358), .A4(new_n752), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND4_X1  g574(.A1(new_n653), .A2(new_n654), .A3(new_n657), .A4(new_n687), .ZN(new_n761));
  INV_X1    g575(.A(new_n752), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n754), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n242), .ZN(G36));
  XNOR2_X1  g578(.A(new_n700), .B(KEYINPUT108), .ZN(new_n765));
  INV_X1    g579(.A(new_n614), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(KEYINPUT43), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n700), .B2(new_n614), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n672), .A2(new_n701), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n520), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n526), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n620), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n739), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n527), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT107), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n785), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n477), .ZN(new_n789));
  INV_X1    g603(.A(new_n751), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n690), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n774), .B2(new_n775), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n776), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  XNOR2_X1  g608(.A(new_n789), .B(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(new_n757), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n796), .A2(new_n722), .A3(new_n238), .A4(new_n751), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n468), .B1(new_n767), .B2(new_n769), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n731), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n710), .A2(new_n711), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT110), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n625), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n802), .B(new_n790), .C1(new_n795), .C2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n800), .B1(new_n807), .B2(KEYINPUT116), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n751), .A2(new_n712), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n734), .ZN(new_n815));
  INV_X1    g629(.A(new_n698), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n238), .A3(new_n469), .A4(new_n809), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n817), .A2(new_n700), .A3(new_n766), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n815), .A2(new_n807), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n712), .A2(new_n600), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT114), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n699), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n802), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n802), .A2(KEYINPUT50), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n808), .B1(new_n819), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n807), .A2(new_n818), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n808), .A2(new_n829), .A3(new_n827), .A4(new_n815), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n615), .ZN(new_n832));
  OAI211_X1 g646(.A(G952), .B(new_n210), .C1(new_n817), .C2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n802), .B2(new_n735), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT48), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n814), .B2(new_n358), .ZN(new_n836));
  AOI211_X1 g650(.A(KEYINPUT48), .B(new_n754), .C1(new_n812), .C2(new_n813), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n834), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n625), .A2(new_n701), .A3(new_n687), .A4(new_n747), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n698), .A2(new_n727), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n688), .A2(new_n706), .A3(new_n736), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT113), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n661), .A2(new_n666), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT101), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n714), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n658), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n603), .B2(new_n604), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n417), .A2(new_n429), .A3(new_n466), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n627), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n681), .A2(new_n862), .A3(new_n724), .A4(new_n732), .ZN(new_n863));
  INV_X1    g677(.A(new_n716), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n615), .A3(new_n627), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n606), .A2(KEYINPUT111), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT111), .B1(new_n606), .B2(new_n865), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n863), .B(new_n864), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n654), .A2(new_n657), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n464), .A2(new_n465), .A3(new_n756), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n625), .A2(new_n679), .A3(new_n624), .A4(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n652), .A3(new_n650), .A4(new_n790), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n331), .A2(new_n336), .B1(G472), .B2(new_n356), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n761), .A2(new_n762), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n875), .B2(new_n358), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n752), .A2(new_n615), .A3(new_n734), .A4(new_n687), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT112), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n757), .A2(new_n879), .A3(new_n734), .A4(new_n752), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n759), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n858), .A2(new_n868), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n854), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n759), .A2(new_n876), .A3(new_n881), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n866), .A2(new_n867), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n863), .A2(new_n864), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n720), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n688), .A2(new_n736), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT52), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n850), .A2(new_n891), .A3(new_n852), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n854), .A2(new_n883), .A3(KEYINPUT53), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n889), .B1(new_n888), .B2(new_n892), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n843), .A2(new_n900), .B1(G952), .B2(G953), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n766), .A2(new_n238), .A3(new_n625), .A4(new_n600), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n699), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n816), .A3(new_n765), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n901), .A2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n210), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(G902), .B1(new_n884), .B2(new_n893), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n911), .B2(G210), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n578), .A2(new_n581), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n579), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n909), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(G902), .C1(new_n884), .C2(new_n893), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n530), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT119), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n916), .B1(new_n924), .B2(new_n926), .ZN(G51));
  XNOR2_X1  g741(.A(new_n894), .B(new_n895), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n739), .B(KEYINPUT57), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n525), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n917), .A2(new_n780), .A3(new_n779), .A4(new_n919), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n908), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND2_X1  g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT120), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n917), .A2(new_n919), .A3(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n647), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n917), .A2(new_n409), .A3(new_n919), .A4(new_n936), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n909), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT121), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n647), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n909), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(G60));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT59), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n928), .A2(new_n612), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n612), .B1(new_n900), .B2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n908), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n894), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n908), .B1(new_n953), .B2(new_n228), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n894), .A2(new_n952), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n955), .A2(KEYINPUT122), .A3(new_n677), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT122), .B1(new_n955), .B2(new_n677), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n954), .B(KEYINPUT61), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  INV_X1    g776(.A(G224), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n472), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n858), .A2(new_n868), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n913), .B1(G898), .B2(new_n210), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT123), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G69));
  AOI21_X1  g783(.A(new_n210), .B1(G227), .B2(G900), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n318), .A2(new_n320), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(new_n400), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(G900), .B2(G953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n763), .B1(new_n795), .B2(new_n797), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n789), .A2(new_n358), .A3(new_n690), .A4(new_n727), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n688), .A2(new_n706), .A3(new_n736), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n759), .A2(new_n974), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n793), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n973), .B1(new_n981), .B2(G953), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n970), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n704), .A2(new_n979), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n692), .A2(new_n751), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n987), .B(new_n358), .C1(new_n615), .C2(new_n861), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n798), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n793), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n972), .B1(new_n992), .B2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n982), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n984), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n984), .A2(new_n994), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n322), .A2(new_n316), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n1000), .B(new_n899), .C1(new_n1001), .C2(new_n342), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n340), .B(KEYINPUT126), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n793), .A2(new_n965), .A3(new_n991), .ZN(new_n1004));
  AOI211_X1 g818(.A(new_n341), .B(new_n1003), .C1(new_n1004), .C2(new_n999), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n341), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n980), .A2(new_n793), .A3(new_n965), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n999), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT127), .B1(new_n1008), .B2(new_n908), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n974), .A2(new_n977), .A3(new_n759), .A4(new_n979), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n776), .B2(new_n792), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1000), .B1(new_n1012), .B2(new_n965), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1010), .B(new_n909), .C1(new_n1013), .C2(new_n1006), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n1002), .B(new_n1005), .C1(new_n1009), .C2(new_n1014), .ZN(G57));
endmodule


