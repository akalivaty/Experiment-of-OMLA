//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G43gat), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n214), .A3(new_n210), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT15), .B1(new_n212), .B2(new_n214), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n209), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n212), .A2(new_n214), .A3(new_n210), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n222), .A2(new_n215), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n209), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n221), .A2(new_n226), .A3(KEYINPUT93), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT93), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n224), .B2(new_n219), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n209), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n202), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  AOI21_X1  g033(.A(G1gat), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(KEYINPUT94), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT95), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(KEYINPUT17), .C1(new_n221), .C2(new_n226), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n221), .A2(new_n226), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT95), .B1(new_n242), .B2(new_n202), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n232), .A2(new_n239), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n239), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n228), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT93), .B1(new_n221), .B2(new_n226), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT96), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n244), .A2(new_n250), .A3(KEYINPUT18), .A4(new_n245), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n245), .B(KEYINPUT13), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n246), .A2(new_n249), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n227), .A2(new_n231), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(new_n239), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT11), .B(G169gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G197gat), .ZN(new_n265));
  XOR2_X1   g064(.A(G113gat), .B(G141gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n251), .A2(KEYINPUT96), .A3(new_n252), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n255), .A2(new_n263), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n268), .B(KEYINPUT91), .ZN(new_n271));
  INV_X1    g070(.A(new_n253), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n262), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G148gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT103), .ZN(new_n279));
  INV_X1    g078(.A(G120gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT102), .ZN(new_n283));
  NAND2_X1  g082(.A1(G85gat), .A2(G92gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT7), .ZN(new_n285));
  NAND2_X1  g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT8), .ZN(new_n287));
  INV_X1    g086(.A(G85gat), .ZN(new_n288));
  INV_X1    g087(.A(G92gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n287), .A2(KEYINPUT98), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT98), .B1(new_n287), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G99gat), .B(G106gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n285), .C1(new_n291), .C2(new_n292), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(KEYINPUT99), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G64gat), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n299), .A2(G57gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(G57gat), .ZN(new_n301));
  AND2_X1   g100(.A1(G71gat), .A2(G78gat), .ZN(new_n302));
  OAI22_X1  g101(.A1(new_n300), .A2(new_n301), .B1(KEYINPUT9), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G71gat), .B(G78gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n291), .A2(new_n292), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT99), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n296), .A4(new_n285), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n298), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n295), .A3(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n283), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  AOI211_X1 g114(.A(KEYINPUT102), .B(new_n313), .C1(new_n310), .C2(new_n311), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT10), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n318), .A3(new_n311), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n309), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT10), .A3(new_n305), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n313), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n282), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT101), .B1(new_n322), .B2(new_n313), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT101), .ZN(new_n326));
  AOI211_X1 g125(.A(new_n326), .B(new_n314), .C1(new_n319), .C2(new_n321), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n317), .B(new_n282), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n328), .B2(KEYINPUT104), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n324), .A2(KEYINPUT104), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(new_n211), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G197gat), .B(G204gat), .Z(new_n336));
  AOI21_X1  g135(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G211gat), .B(G218gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT74), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n338), .A2(KEYINPUT74), .A3(new_n339), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(new_n347), .B2(KEYINPUT77), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n349), .B(new_n350), .C1(G155gat), .C2(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G141gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G148gat), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G141gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n354), .A2(new_n356), .B1(KEYINPUT2), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(G155gat), .B(G162gat), .C1(new_n352), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(KEYINPUT2), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(new_n357), .A3(new_n348), .A4(new_n351), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n347), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n359), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n346), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n345), .A2(new_n367), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n364), .ZN(new_n373));
  OAI211_X1 g172(.A(G228gat), .B(G233gat), .C1(new_n370), .C2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n340), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n367), .B1(new_n377), .B2(new_n342), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(KEYINPUT85), .B2(new_n342), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n369), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n335), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(G22gat), .Z(new_n386));
  NAND3_X1  g185(.A1(new_n374), .A2(new_n335), .A3(new_n382), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n384), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  INV_X1    g190(.A(G183gat), .ZN(new_n392));
  INV_X1    g191(.A(G190gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n394), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT23), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n400), .B(new_n405), .C1(new_n406), .C2(new_n402), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT25), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n401), .B1(KEYINPUT23), .B2(new_n403), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n397), .A2(new_n398), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n393), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT64), .B(G169gat), .Z(new_n413));
  NOR2_X1   g212(.A1(new_n406), .A2(G176gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT25), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT27), .B1(new_n392), .B2(KEYINPUT66), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT27), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G183gat), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n418), .B(new_n393), .C1(KEYINPUT66), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT28), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT27), .B(G183gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(G190gat), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n395), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n402), .A2(KEYINPUT26), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT26), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n427), .A2(new_n403), .A3(new_n429), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT70), .B1(new_n417), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G127gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(G134gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT67), .B(G127gat), .ZN(new_n436));
  INV_X1    g235(.A(G134gat), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT68), .B(new_n435), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT67), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(G127gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n433), .A2(KEYINPUT67), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n439), .B(G134gat), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G113gat), .B(G120gat), .Z(new_n444));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n438), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n437), .A2(G127gat), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n434), .A2(new_n450), .A3(KEYINPUT1), .ZN(new_n451));
  XNOR2_X1  g250(.A(G113gat), .B(G120gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT69), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n407), .A2(KEYINPUT25), .B1(new_n412), .B2(new_n415), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n427), .A2(new_n403), .A3(new_n429), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n392), .A2(KEYINPUT27), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n460));
  AOI21_X1  g259(.A(G190gat), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT28), .B1(new_n461), .B2(new_n418), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n423), .A2(new_n424), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n395), .B(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n432), .A2(new_n455), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G227gat), .ZN(new_n467));
  INV_X1    g266(.A(G233gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n456), .A2(new_n464), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n447), .A2(new_n454), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT32), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT72), .B(G71gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G99gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT71), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n473), .A2(new_n482), .A3(KEYINPUT32), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n475), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT73), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n485), .B2(new_n479), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(KEYINPUT32), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT34), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n466), .A2(new_n472), .ZN(new_n491));
  INV_X1    g290(.A(new_n469), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n484), .A2(new_n495), .A3(new_n488), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n495), .B1(new_n484), .B2(new_n488), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n390), .A2(KEYINPUT35), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n371), .A2(new_n471), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT4), .B1(new_n375), .B2(new_n455), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT79), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n447), .A2(new_n508), .A3(new_n454), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n447), .B2(new_n454), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n366), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n375), .A2(new_n455), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT80), .A3(new_n502), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n506), .A2(new_n512), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n513), .ZN(new_n517));
  INV_X1    g316(.A(new_n511), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n371), .B1(new_n518), .B2(new_n509), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n519), .B2(new_n514), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(KEYINPUT5), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT81), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT81), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n516), .A2(new_n523), .A3(KEYINPUT5), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT83), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT83), .B1(new_n503), .B2(new_n504), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT5), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n530), .A3(new_n513), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G1gat), .B(G29gat), .Z(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G85gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(KEYINPUT6), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n539), .A3(new_n533), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n532), .B1(new_n522), .B2(new_n524), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G226gat), .A2(G233gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n417), .A2(new_n431), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(KEYINPUT29), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT75), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n548), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n470), .A2(new_n367), .B1(G226gat), .B2(G233gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n551), .B(new_n346), .C1(new_n554), .C2(KEYINPUT75), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n345), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G36gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(new_n236), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT30), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n555), .B2(new_n556), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI211_X1 g364(.A(KEYINPUT30), .B(new_n561), .C1(new_n555), .C2(new_n556), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n547), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n501), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n498), .A2(new_n493), .A3(new_n499), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n494), .B1(new_n490), .B2(new_n496), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT6), .B1(new_n545), .B2(new_n539), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n540), .B1(new_n545), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g375(.A(KEYINPUT88), .B(new_n532), .C1(new_n522), .C2(new_n524), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n541), .A2(KEYINPUT90), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT90), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n546), .A2(new_n580), .A3(KEYINPUT6), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n573), .A2(new_n582), .A3(new_n567), .A4(new_n390), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n569), .B1(new_n570), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n571), .B2(new_n572), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n500), .A2(new_n497), .A3(KEYINPUT36), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n388), .A2(new_n389), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n586), .A2(new_n587), .B1(new_n568), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n512), .ZN(new_n590));
  INV_X1    g389(.A(new_n528), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(new_n526), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT86), .B1(new_n592), .B2(new_n513), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT86), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(new_n517), .C1(new_n529), .C2(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OR3_X1    g397(.A1(new_n519), .A2(new_n517), .A3(new_n514), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT39), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n600), .A3(new_n539), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n545), .A2(new_n575), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n540), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n565), .A2(new_n566), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n598), .A2(new_n600), .A3(KEYINPUT40), .A4(new_n539), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n562), .B1(new_n557), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n555), .A2(KEYINPUT37), .A3(new_n556), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n564), .B1(new_n613), .B2(KEYINPUT38), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n578), .A2(new_n579), .A3(new_n614), .A4(new_n581), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n554), .A2(new_n345), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT89), .Z(new_n617));
  OAI211_X1 g416(.A(new_n345), .B(new_n551), .C1(new_n554), .C2(KEYINPUT75), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT37), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n620), .A2(new_n621), .A3(new_n611), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n390), .B(new_n609), .C1(new_n615), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n589), .A2(new_n623), .ZN(new_n624));
  AOI211_X1 g423(.A(new_n276), .B(new_n332), .C1(new_n584), .C2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT21), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n239), .B1(new_n626), .B2(new_n306), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G183gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n305), .A2(KEYINPUT21), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n633), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n320), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n232), .A2(new_n639), .A3(new_n241), .A4(new_n243), .ZN(new_n640));
  NAND2_X1  g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n249), .B2(new_n320), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT100), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G134gat), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n641), .A2(new_n642), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT97), .ZN(new_n651));
  INV_X1    g450(.A(G162gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n648), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n649), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n649), .B2(new_n654), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n625), .A2(new_n638), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n547), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g462(.A1(new_n659), .A2(new_n567), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n234), .A2(new_n236), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(new_n669), .C1(new_n236), .C2(new_n664), .ZN(G1325gat));
  NAND2_X1  g469(.A1(new_n586), .A2(new_n587), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n660), .A2(G15gat), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n573), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(G15gat), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT105), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n659), .A2(new_n390), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT106), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n678), .B(new_n680), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n638), .A2(new_n658), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n625), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n203), .A3(new_n661), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n331), .B(KEYINPUT107), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n276), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n657), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n624), .A2(KEYINPUT108), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n589), .A2(new_n623), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n584), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT109), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n690), .A2(new_n695), .A3(new_n584), .A4(new_n692), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n689), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n584), .A2(new_n624), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n688), .B1(new_n698), .B2(new_n657), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n637), .B(new_n687), .C1(new_n697), .C2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n547), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n701), .ZN(G1328gat));
  OAI21_X1  g501(.A(G36gat), .B1(new_n700), .B2(new_n567), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n204), .A3(new_n607), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(KEYINPUT110), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n705), .A2(KEYINPUT110), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n703), .B(new_n708), .C1(new_n706), .C2(new_n704), .ZN(G1329gat));
  NOR3_X1   g508(.A1(new_n700), .A2(new_n213), .A3(new_n671), .ZN(new_n710));
  AOI21_X1  g509(.A(G43gat), .B1(new_n683), .B2(new_n573), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n710), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT47), .B1(new_n710), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n700), .B2(new_n390), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n683), .A2(new_n211), .A3(new_n588), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1331gat));
  INV_X1    g518(.A(new_n686), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n694), .B2(new_n696), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n637), .A2(new_n657), .A3(new_n275), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n661), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n567), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  NAND3_X1  g530(.A1(new_n724), .A2(G71gat), .A3(new_n672), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n723), .A2(new_n674), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(G71gat), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n723), .A2(new_n390), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT111), .B(G78gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1335gat));
  NAND3_X1  g537(.A1(new_n693), .A2(new_n276), .A3(new_n682), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT51), .Z(new_n740));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n547), .A2(G85gat), .A3(new_n331), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT113), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n637), .B(new_n276), .C1(new_n697), .C2(new_n699), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n746), .A2(new_n547), .A3(new_n331), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n288), .B2(new_n747), .ZN(G1336gat));
  NAND4_X1  g547(.A1(new_n740), .A2(new_n289), .A3(new_n607), .A4(new_n686), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n746), .A2(new_n567), .A3(new_n331), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n289), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n753), .B(new_n749), .C1(new_n750), .C2(new_n289), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1337gat));
  NOR3_X1   g554(.A1(new_n674), .A2(new_n331), .A3(G99gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n742), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G99gat), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n746), .A2(new_n671), .A3(new_n331), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(G1338gat));
  INV_X1    g559(.A(G106gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n761), .A3(new_n588), .A4(new_n686), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n390), .A3(new_n331), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n761), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT53), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n766), .B(new_n762), .C1(new_n763), .C2(new_n761), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1339gat));
  NOR4_X1   g567(.A1(new_n637), .A2(new_n657), .A3(new_n275), .A4(new_n332), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n260), .A2(new_n239), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n250), .A2(new_n770), .A3(new_n257), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT116), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n245), .B1(new_n244), .B2(new_n250), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n267), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n657), .A2(new_n270), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n328), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n281), .B1(new_n323), .B2(KEYINPUT54), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n323), .A2(new_n326), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n314), .B1(new_n319), .B2(new_n321), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT101), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n319), .A2(new_n314), .A3(new_n321), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n778), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n777), .B1(new_n785), .B2(KEYINPUT55), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n325), .B2(new_n327), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n282), .B1(new_n780), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g592(.A(KEYINPUT114), .B(KEYINPUT55), .C1(new_n788), .C2(new_n790), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n786), .B(new_n797), .C1(new_n793), .C2(new_n794), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n776), .A2(new_n796), .A3(KEYINPUT117), .A4(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n796), .A2(new_n275), .A3(new_n798), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n774), .B(new_n270), .C1(new_n329), .C2(new_n330), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(KEYINPUT118), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n658), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT118), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n769), .B1(new_n809), .B2(new_n637), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n674), .A2(new_n588), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n661), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n607), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(KEYINPUT119), .A3(new_n661), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n276), .A2(G113gat), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT120), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n813), .A2(new_n661), .A3(new_n567), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n276), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1340gat));
  NAND3_X1  g623(.A1(new_n818), .A2(new_n280), .A3(new_n332), .ZN(new_n825));
  OAI21_X1  g624(.A(G120gat), .B1(new_n822), .B2(new_n720), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1341gat));
  INV_X1    g626(.A(new_n436), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n822), .A2(new_n828), .A3(new_n637), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n818), .A2(new_n638), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n828), .ZN(G1342gat));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n437), .A3(new_n657), .A4(new_n817), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n822), .B2(new_n658), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  NAND2_X1  g635(.A1(new_n804), .A2(new_n805), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n658), .A3(new_n806), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n638), .B1(new_n840), .B2(new_n803), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n588), .B1(new_n841), .B2(new_n769), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n661), .A2(new_n567), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n672), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n353), .A3(new_n275), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n791), .A2(new_n792), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n275), .A2(new_n786), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n805), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n852), .A3(new_n805), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n658), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n638), .B1(new_n803), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n588), .B1(new_n855), .B2(new_n769), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT57), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n844), .B(new_n857), .C1(new_n842), .C2(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n276), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n847), .B1(new_n859), .B2(new_n353), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT58), .ZN(G1344gat));
  OR2_X1    g660(.A1(new_n775), .A2(new_n795), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n854), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n854), .A2(KEYINPUT123), .A3(new_n862), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n637), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n769), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n842), .A2(KEYINPUT57), .B1(new_n869), .B2(new_n588), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  AOI211_X1 g670(.A(new_n871), .B(new_n331), .C1(new_n845), .C2(KEYINPUT122), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n870), .B(new_n872), .C1(KEYINPUT122), .C2(new_n845), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n858), .B2(new_n331), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n355), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(G148gat), .B1(new_n846), .B2(new_n332), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(KEYINPUT59), .B2(new_n876), .ZN(G1345gat));
  AOI21_X1  g676(.A(G155gat), .B1(new_n846), .B2(new_n638), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n858), .A2(new_n637), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n846), .B2(new_n657), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n858), .A2(new_n652), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n657), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n661), .A2(new_n567), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n813), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n413), .A3(new_n275), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(KEYINPUT124), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n813), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n276), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G169gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n886), .B2(new_n332), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n888), .A2(new_n890), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(G176gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(new_n686), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n886), .A2(new_n638), .A3(new_n423), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n637), .B1(new_n888), .B2(new_n890), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n392), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n902), .B(new_n898), .C1(new_n899), .C2(new_n392), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n393), .A3(new_n657), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n895), .A2(new_n657), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(G190gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n658), .B1(new_n888), .B2(new_n890), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(KEYINPUT61), .A3(new_n393), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n908), .B2(new_n910), .ZN(G1351gat));
  AND2_X1   g710(.A1(new_n671), .A2(new_n884), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n870), .A2(new_n275), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G197gat), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n588), .B(new_n912), .C1(new_n841), .C2(new_n769), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n276), .A2(G197gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(G1352gat));
  NAND3_X1  g716(.A1(new_n870), .A2(new_n686), .A3(new_n912), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G204gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n915), .A2(G204gat), .A3(new_n331), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(G1353gat));
  OAI21_X1  g723(.A(KEYINPUT57), .B1(new_n810), .B2(new_n390), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n854), .A2(KEYINPUT123), .A3(new_n862), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT123), .B1(new_n854), .B2(new_n862), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(new_n638), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n926), .B(new_n588), .C1(new_n929), .C2(new_n769), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n925), .A2(new_n638), .A3(new_n930), .A4(new_n912), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n933), .A2(G211gat), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  OR3_X1    g738(.A1(new_n915), .A2(G211gat), .A3(new_n637), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n870), .A2(new_n932), .A3(new_n638), .A4(new_n912), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n931), .A2(KEYINPUT125), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n941), .A2(new_n942), .A3(G211gat), .A4(new_n938), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n936), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n939), .A2(new_n940), .A3(new_n944), .ZN(G1354gat));
  NAND3_X1  g744(.A1(new_n870), .A2(new_n657), .A3(new_n912), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G218gat), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n658), .A2(G218gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n915), .B2(new_n948), .ZN(G1355gat));
endmodule


