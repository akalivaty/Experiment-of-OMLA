//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n462), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n462), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n467), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n473), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(G162));
  NOR2_X1   g058(.A1(new_n462), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n479), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n462), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .A3(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n486), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n463), .A2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n462), .A3(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n499), .A2(new_n462), .A3(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n467), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n496), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI211_X1 g083(.A(KEYINPUT72), .B(new_n507), .C1(new_n508), .C2(KEYINPUT73), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT5), .B1(new_n508), .B2(KEYINPUT72), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(new_n519), .B1(KEYINPUT6), .B2(new_n515), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n515), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(new_n514), .A2(new_n520), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n520), .A2(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n530), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n521), .A2(new_n541), .B1(new_n523), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n515), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n521), .A2(new_n547), .B1(new_n523), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n559), .A2(new_n560), .B1(G91), .B2(new_n529), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n514), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G65), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n515), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  OR2_X1    g146(.A1(G166), .A2(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g147(.A1(G166), .A2(KEYINPUT78), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(G303));
  NAND2_X1  g149(.A1(new_n529), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n531), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n514), .A2(G61), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(new_n580), .B1(G73), .B2(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n514), .A2(KEYINPUT79), .A3(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n521), .A2(new_n585), .B1(new_n523), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  AND2_X1   g164(.A1(new_n514), .A2(G60), .ZN(new_n590));
  AND2_X1   g165(.A1(G72), .A2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  AOI22_X1  g170(.A1(G85), .A2(new_n529), .B1(new_n531), .B2(G47), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n564), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n515), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(new_n599), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n521), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n603), .A2(new_n606), .B1(G54), .B2(new_n531), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT82), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n568), .A2(KEYINPUT83), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n568), .A2(KEYINPUT83), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(G297));
  XOR2_X1   g193(.A(G297), .B(KEYINPUT84), .Z(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n609), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND3_X1  g196(.A1(new_n602), .A2(new_n620), .A3(new_n607), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n492), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n462), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G135), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n626), .B1(new_n627), .B2(new_n628), .C1(new_n629), .C2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n467), .A2(new_n471), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n631), .B1(G2100), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(G2100), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(KEYINPUT86), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(KEYINPUT86), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT87), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n647), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT88), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT89), .ZN(new_n660));
  NOR2_X1   g235(.A1(G2072), .A2(G2078), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n442), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(new_n662), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n662), .B(KEYINPUT17), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n664), .C1(new_n660), .C2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n660), .A2(new_n668), .A3(new_n663), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n686), .B(new_n685), .S(new_n678), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1981), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(G1986), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(G1986), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n689), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n694), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n675), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n694), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(new_n702), .A3(new_n674), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(G229));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT92), .B1(G95), .B2(G2105), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g284(.A1(KEYINPUT92), .A2(G95), .A3(G2105), .ZN(new_n710));
  OAI221_X1 g285(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n492), .A2(G119), .ZN(new_n712));
  INV_X1    g287(.A(G131), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n473), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT91), .B(G29), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G25), .B(new_n714), .S(new_n716), .Z(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT35), .B(G1991), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n587), .B1(new_n583), .B2(G651), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G6), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT32), .B(G1981), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G22), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G166), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(G23), .ZN(new_n732));
  INV_X1    g307(.A(G288), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n727), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT33), .B(G1976), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n725), .A2(new_n726), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n719), .B1(new_n737), .B2(KEYINPUT34), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n707), .B(new_n738), .C1(KEYINPUT34), .C2(new_n737), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT36), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G139), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n473), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  INV_X1    g323(.A(G127), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n497), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n747), .B1(G2105), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT95), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n742), .B1(new_n752), .B2(new_n741), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G2072), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n715), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n482), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n492), .A2(G128), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n741), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G29), .B2(G32), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n492), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n741), .ZN(new_n773));
  MUX2_X1   g348(.A(new_n767), .B(new_n766), .S(new_n773), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n765), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n727), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  INV_X1    g356(.A(G19), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n782), .A2(KEYINPUT94), .A3(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(KEYINPUT94), .B1(new_n782), .B2(G16), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n783), .B(new_n784), .C1(new_n552), .C2(new_n727), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n754), .A2(new_n777), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n609), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G4), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT30), .B(G28), .ZN(new_n792));
  OR2_X1    g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  NAND2_X1  g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n792), .A2(new_n741), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n630), .B2(new_n715), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n716), .A2(G35), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n716), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT98), .B(G2090), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n798), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G164), .A2(new_n715), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G27), .B2(new_n715), .ZN(new_n804));
  INV_X1    g379(.A(G2078), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n796), .B(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n727), .A2(G5), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G171), .B2(new_n727), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT24), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(G34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(G34), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n715), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G160), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n741), .ZN(new_n815));
  INV_X1    g390(.A(G2084), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n809), .A2(G1961), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n809), .A2(G1961), .B1(new_n815), .B2(new_n816), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n806), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n727), .A2(G21), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G168), .B2(new_n727), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1966), .ZN(new_n823));
  NOR4_X1   g398(.A1(new_n787), .A2(new_n791), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n740), .A2(KEYINPUT99), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT99), .B1(new_n740), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n740), .A2(new_n824), .ZN(G150));
  NAND2_X1  g403(.A1(new_n609), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT101), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(G93), .A2(new_n529), .B1(new_n531), .B2(G55), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n515), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n552), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n832), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT102), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  OR2_X1    g418(.A1(new_n840), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(G160), .B(new_n630), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  INV_X1    g421(.A(new_n772), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n752), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n752), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n492), .A2(G130), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT104), .Z(new_n851));
  INV_X1    g426(.A(G118), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(KEYINPUT105), .A3(G2105), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT105), .B1(new_n852), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n482), .A2(G142), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n714), .ZN(new_n859));
  OR3_X1    g434(.A1(new_n848), .A2(new_n849), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n848), .B2(new_n849), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR4_X1   g437(.A1(new_n497), .A2(new_n487), .A3(new_n488), .A4(new_n462), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT69), .B1(new_n492), .B2(G126), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n863), .A2(new_n864), .B1(new_n484), .B2(new_n485), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n504), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n498), .B1(new_n497), .B2(new_n500), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n467), .A2(new_n502), .A3(KEYINPUT70), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(KEYINPUT103), .A3(new_n496), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n865), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n761), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n634), .Z(new_n874));
  NOR2_X1   g449(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n860), .A2(new_n861), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n846), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n862), .A2(new_n874), .ZN(new_n881));
  INV_X1    g456(.A(new_n846), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g461(.A(KEYINPUT106), .B1(new_n835), .B2(new_n615), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n622), .A2(new_n836), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n622), .A2(new_n836), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n602), .A2(new_n568), .A3(new_n607), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n568), .B1(new_n602), .B2(new_n607), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n892), .B2(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(new_n893), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n890), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n897), .A2(new_n899), .B1(new_n888), .B2(new_n889), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n890), .A2(new_n894), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G290), .B(G305), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n733), .B(G166), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n907), .B(new_n908), .Z(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G868), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n903), .B2(new_n906), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n887), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n915), .A2(KEYINPUT106), .A3(G868), .A4(new_n911), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(G295));
  AND3_X1   g492(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT107), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT107), .B1(new_n914), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(G331));
  XNOR2_X1  g495(.A(G168), .B(G301), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n836), .ZN(new_n922));
  INV_X1    g497(.A(new_n836), .ZN(new_n923));
  NOR2_X1   g498(.A1(G286), .A2(G301), .ZN(new_n924));
  NOR2_X1   g499(.A1(G168), .A2(G171), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n897), .A3(new_n899), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n926), .A3(new_n894), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n909), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n910), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n880), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n935), .A3(new_n880), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(G397));
  AOI221_X4 g514(.A(new_n866), .B1(new_n495), .B2(KEYINPUT4), .C1(new_n868), .C2(new_n869), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT103), .B1(new_n870), .B2(new_n496), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n494), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT45), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n475), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n466), .A2(new_n469), .ZN(new_n947));
  OAI211_X1 g522(.A(G40), .B(new_n946), .C1(new_n947), .C2(new_n462), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1996), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n772), .B(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n761), .B(new_n764), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n714), .B(new_n718), .Z(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n942), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n505), .A2(new_n943), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n470), .A2(new_n964), .A3(new_n475), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n730), .ZN(new_n967));
  INV_X1    g542(.A(G2090), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT50), .B1(new_n942), .B2(new_n943), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n494), .B2(new_n504), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n968), .B(new_n965), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT108), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n572), .A2(G8), .A3(new_n573), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(KEYINPUT55), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n976), .A2(KEYINPUT55), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n975), .B1(new_n979), .B2(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n967), .A2(new_n982), .A3(new_n972), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n974), .A2(new_n981), .A3(G8), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n967), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n948), .B1(new_n970), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n872), .A2(G1384), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(new_n986), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(G2090), .ZN(new_n990));
  OAI21_X1  g565(.A(G8), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n980), .A3(new_n978), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n948), .A2(G2084), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n969), .B2(new_n971), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT115), .ZN(new_n996));
  INV_X1    g571(.A(G1966), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n965), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n944), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n994), .C1(new_n969), .C2(new_n971), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n996), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(G8), .A3(G168), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G305), .A2(G1981), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(new_n720), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n515), .B1(new_n581), .B2(new_n582), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n1010), .A2(KEYINPUT112), .A3(G1981), .A4(new_n587), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n872), .A2(new_n948), .A3(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT110), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n942), .A2(new_n943), .A3(new_n965), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(G8), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1012), .A2(new_n1013), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n720), .A2(new_n1008), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(G305), .B2(G1981), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1011), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n733), .A2(G1976), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1017), .A2(new_n1018), .A3(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1018), .B1(new_n1017), .B2(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1020), .A2(new_n1025), .B1(new_n1029), .B2(KEYINPUT52), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1026), .B(new_n1032), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1026), .A4(new_n1032), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1030), .A2(new_n1038), .A3(KEYINPUT114), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT114), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n993), .B(new_n1005), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1005), .A2(new_n984), .A3(KEYINPUT63), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n974), .A2(G8), .A3(new_n983), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n980), .A3(new_n978), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1044), .A2(new_n1038), .A3(new_n1030), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n996), .A2(G168), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1015), .A2(KEYINPUT120), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1003), .A2(G8), .A3(G286), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1052), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1050), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1057), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(KEYINPUT62), .A3(new_n1055), .A4(new_n1054), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n960), .A2(new_n963), .A3(new_n805), .A4(new_n965), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(KEYINPUT121), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT121), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n965), .B1(new_n969), .B2(new_n971), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1063), .A2(G2078), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n945), .A2(new_n965), .A3(new_n1070), .A4(new_n998), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(G171), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n993), .B(new_n1074), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1049), .B1(new_n1061), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n733), .A2(new_n1031), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1035), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1030), .A2(new_n1038), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n984), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT113), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n984), .A2(new_n992), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1035), .B1(new_n1024), .B2(KEYINPUT49), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1085), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1030), .A2(new_n1038), .A3(KEYINPUT114), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1084), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(KEYINPUT124), .A4(new_n1074), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1048), .A2(new_n1076), .A3(new_n1083), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1056), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1065), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1062), .A2(KEYINPUT121), .A3(new_n1063), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1072), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1101), .B2(G301), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n948), .B1(new_n988), .B2(KEYINPUT45), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n945), .A3(new_n1070), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(KEYINPUT122), .A3(new_n945), .A4(new_n1070), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1069), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(G171), .B1(new_n1108), .B2(new_n1066), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1097), .A2(new_n1059), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1107), .A2(new_n1069), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(G301), .A4(new_n1106), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1073), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1111), .B1(new_n1115), .B2(new_n1098), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1114), .C2(new_n1073), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1093), .B(new_n1110), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n565), .A2(new_n566), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1119), .B(new_n561), .C1(new_n1120), .C2(new_n515), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT57), .B1(new_n562), .B2(new_n567), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1103), .A2(new_n963), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1956), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n989), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1067), .A2(new_n790), .B1(new_n764), .B2(new_n1014), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n608), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1128), .B1(new_n1131), .B2(KEYINPUT116), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(KEYINPUT116), .B2(new_n1131), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1125), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1125), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT61), .B1(new_n1136), .B2(new_n1128), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1123), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1134), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n960), .A2(new_n963), .A3(new_n950), .A4(new_n965), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  AND3_X1   g721(.A1(new_n1017), .A2(KEYINPUT117), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT117), .B1(new_n1017), .B2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT118), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(new_n1145), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1144), .B1(new_n1153), .B2(new_n552), .ZN(new_n1154));
  INV_X1    g729(.A(new_n552), .ZN(new_n1155));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n1155), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1143), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1143), .B(KEYINPUT119), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(new_n609), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(KEYINPUT60), .B2(new_n1129), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1118), .B1(new_n1135), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n959), .B1(new_n1096), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n955), .A2(new_n949), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n949), .A2(new_n956), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT126), .Z(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1169), .B2(KEYINPUT48), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(KEYINPUT48), .B2(new_n1169), .ZN(new_n1171));
  INV_X1    g746(.A(new_n949), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1172), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT46), .B1(new_n1172), .B2(G1996), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n952), .A2(new_n847), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1174), .B1(new_n949), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT47), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n714), .A2(new_n718), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1172), .B2(new_n953), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(G2067), .B2(new_n761), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n949), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1171), .A2(new_n1177), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1166), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(G319), .ZN(new_n1187));
  NOR2_X1   g761(.A1(G227), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n657), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n700), .B2(new_n703), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1190), .A2(new_n885), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1191), .B1(new_n934), .B2(new_n936), .ZN(new_n1192));
  XNOR2_X1  g766(.A(new_n1192), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g767(.A(new_n1192), .ZN(G225));
endmodule


