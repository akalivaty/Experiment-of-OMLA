

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n582, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723;

  XNOR2_X1 U368 ( .A(KEYINPUT32), .B(n573), .ZN(n722) );
  NOR2_X1 U369 ( .A1(n639), .A2(n640), .ZN(n636) );
  AND2_X1 U370 ( .A1(n395), .A2(n393), .ZN(n392) );
  XNOR2_X1 U371 ( .A(n708), .B(G146), .ZN(n477) );
  XOR2_X1 U372 ( .A(G137), .B(G140), .Z(n454) );
  NOR2_X2 U373 ( .A1(n392), .A2(n388), .ZN(n387) );
  XNOR2_X1 U374 ( .A(n346), .B(n353), .ZN(n381) );
  NAND2_X1 U375 ( .A1(n672), .A2(n580), .ZN(n346) );
  NAND2_X1 U376 ( .A1(n347), .A2(n584), .ZN(n601) );
  XNOR2_X1 U377 ( .A(n398), .B(n397), .ZN(n347) );
  NAND2_X1 U378 ( .A1(n636), .A2(n542), .ZN(n470) );
  NOR2_X2 U379 ( .A1(n687), .A2(n696), .ZN(n367) );
  NAND2_X2 U380 ( .A1(n633), .A2(n602), .ZN(n604) );
  OR2_X2 U381 ( .A1(n678), .A2(n602), .ZN(n382) );
  NAND2_X1 U382 ( .A1(n616), .A2(n722), .ZN(n596) );
  AND2_X1 U383 ( .A1(n637), .A2(n636), .ZN(n588) );
  AND2_X1 U384 ( .A1(n357), .A2(n354), .ZN(n379) );
  NOR2_X1 U385 ( .A1(n551), .A2(n550), .ZN(n654) );
  XNOR2_X1 U386 ( .A(n468), .B(KEYINPUT68), .ZN(n469) );
  INV_X4 U387 ( .A(G953), .ZN(n455) );
  AND2_X2 U388 ( .A1(n360), .A2(n359), .ZN(n603) );
  XNOR2_X2 U389 ( .A(n513), .B(n433), .ZN(n708) );
  XNOR2_X1 U390 ( .A(n456), .B(n457), .ZN(n514) );
  NOR2_X1 U391 ( .A1(n400), .A2(n656), .ZN(n539) );
  XNOR2_X1 U392 ( .A(G131), .B(KEYINPUT4), .ZN(n433) );
  AND2_X1 U393 ( .A1(n416), .A2(n415), .ZN(n599) );
  INV_X1 U394 ( .A(KEYINPUT65), .ZN(n397) );
  NOR2_X1 U395 ( .A1(n361), .A2(KEYINPUT44), .ZN(n398) );
  XNOR2_X1 U396 ( .A(G143), .B(G140), .ZN(n501) );
  NOR2_X1 U397 ( .A1(n622), .A2(n545), .ZN(n557) );
  NAND2_X1 U398 ( .A1(n391), .A2(n390), .ZN(n389) );
  AND2_X1 U399 ( .A1(n469), .A2(n394), .ZN(n390) );
  INV_X1 U400 ( .A(KEYINPUT1), .ZN(n388) );
  AND2_X1 U401 ( .A1(n389), .A2(n388), .ZN(n385) );
  OR2_X1 U402 ( .A1(n469), .A2(n394), .ZN(n393) );
  INV_X1 U403 ( .A(n469), .ZN(n396) );
  XNOR2_X1 U404 ( .A(n481), .B(n480), .ZN(n543) );
  XNOR2_X1 U405 ( .A(G101), .B(G137), .ZN(n473) );
  XOR2_X1 U406 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n474) );
  XNOR2_X1 U407 ( .A(n351), .B(n443), .ZN(n478) );
  XNOR2_X1 U408 ( .A(KEYINPUT3), .B(G119), .ZN(n443) );
  INV_X1 U409 ( .A(KEYINPUT24), .ZN(n459) );
  XNOR2_X1 U410 ( .A(G119), .B(G110), .ZN(n460) );
  XOR2_X1 U411 ( .A(G128), .B(KEYINPUT23), .Z(n458) );
  XNOR2_X1 U412 ( .A(G107), .B(G122), .ZN(n518) );
  INV_X1 U413 ( .A(KEYINPUT9), .ZN(n376) );
  XOR2_X1 U414 ( .A(G116), .B(KEYINPUT7), .Z(n516) );
  XOR2_X1 U415 ( .A(G146), .B(G125), .Z(n453) );
  XNOR2_X1 U416 ( .A(n441), .B(n426), .ZN(n425) );
  XNOR2_X1 U417 ( .A(KEYINPUT17), .B(KEYINPUT72), .ZN(n426) );
  XNOR2_X1 U418 ( .A(n424), .B(KEYINPUT18), .ZN(n423) );
  XNOR2_X1 U419 ( .A(KEYINPUT4), .B(KEYINPUT86), .ZN(n424) );
  NOR2_X1 U420 ( .A1(n653), .A2(n552), .ZN(n492) );
  XNOR2_X1 U421 ( .A(n371), .B(n355), .ZN(n574) );
  NOR2_X1 U422 ( .A1(n591), .A2(n421), .ZN(n371) );
  NAND2_X1 U423 ( .A1(n654), .A2(n526), .ZN(n421) );
  XNOR2_X1 U424 ( .A(n547), .B(KEYINPUT19), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n464), .B(n365), .ZN(n413) );
  XNOR2_X1 U426 ( .A(n466), .B(KEYINPUT25), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n362), .B(n444), .ZN(n697) );
  XNOR2_X1 U428 ( .A(n478), .B(n445), .ZN(n362) );
  XOR2_X1 U429 ( .A(G122), .B(KEYINPUT16), .Z(n445) );
  INV_X1 U430 ( .A(G902), .ZN(n394) );
  OR2_X1 U431 ( .A1(G237), .A2(G902), .ZN(n471) );
  NAND2_X1 U432 ( .A1(n549), .A2(n556), .ZN(n409) );
  OR2_X1 U433 ( .A1(n720), .A2(n412), .ZN(n408) );
  INV_X1 U434 ( .A(n630), .ZN(n410) );
  NAND2_X1 U435 ( .A1(n554), .A2(n411), .ZN(n406) );
  XNOR2_X1 U436 ( .A(n440), .B(KEYINPUT85), .ZN(n602) );
  XNOR2_X1 U437 ( .A(G902), .B(KEYINPUT15), .ZN(n440) );
  NAND2_X1 U438 ( .A1(n414), .A2(n640), .ZN(n528) );
  AND2_X1 U439 ( .A1(n526), .A2(n527), .ZN(n414) );
  XNOR2_X1 U440 ( .A(n377), .B(KEYINPUT45), .ZN(n360) );
  NAND2_X1 U441 ( .A1(n600), .A2(n601), .ZN(n377) );
  XNOR2_X1 U442 ( .A(G113), .B(G131), .ZN(n499) );
  NOR2_X1 U443 ( .A1(n389), .A2(n388), .ZN(n386) );
  NOR2_X1 U444 ( .A1(n592), .A2(n483), .ZN(n490) );
  INV_X1 U445 ( .A(KEYINPUT0), .ZN(n422) );
  XNOR2_X1 U446 ( .A(n476), .B(n374), .ZN(n373) );
  XNOR2_X1 U447 ( .A(n402), .B(n401), .ZN(n462) );
  XNOR2_X1 U448 ( .A(n461), .B(n458), .ZN(n402) );
  NAND2_X1 U449 ( .A1(n514), .A2(G221), .ZN(n401) );
  XNOR2_X1 U450 ( .A(n517), .B(n375), .ZN(n519) );
  XNOR2_X1 U451 ( .A(n518), .B(n376), .ZN(n375) );
  NAND2_X1 U452 ( .A1(n688), .A2(G469), .ZN(n420) );
  XNOR2_X1 U453 ( .A(n363), .B(n697), .ZN(n678) );
  XNOR2_X1 U454 ( .A(n425), .B(n423), .ZN(n442) );
  INV_X1 U455 ( .A(n582), .ZN(n380) );
  XNOR2_X1 U456 ( .A(n537), .B(KEYINPUT74), .ZN(n400) );
  INV_X1 U457 ( .A(n536), .ZN(n358) );
  INV_X1 U458 ( .A(KEYINPUT53), .ZN(n369) );
  AND2_X1 U459 ( .A1(n637), .A2(n372), .ZN(n348) );
  NOR2_X1 U460 ( .A1(n669), .A2(G953), .ZN(n349) );
  XOR2_X1 U461 ( .A(G104), .B(G107), .Z(n350) );
  XOR2_X1 U462 ( .A(G113), .B(G116), .Z(n351) );
  NOR2_X1 U463 ( .A1(n720), .A2(n406), .ZN(n352) );
  XNOR2_X1 U464 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n353) );
  OR2_X1 U465 ( .A1(n571), .A2(n570), .ZN(n354) );
  XOR2_X1 U466 ( .A(KEYINPUT22), .B(KEYINPUT71), .Z(n355) );
  XNOR2_X1 U467 ( .A(n477), .B(n373), .ZN(n606) );
  XOR2_X1 U468 ( .A(n606), .B(KEYINPUT62), .Z(n356) );
  NOR2_X1 U469 ( .A1(G952), .A2(n455), .ZN(n696) );
  INV_X1 U470 ( .A(n696), .ZN(n418) );
  NAND2_X1 U471 ( .A1(n358), .A2(n357), .ZN(n537) );
  INV_X1 U472 ( .A(n713), .ZN(n359) );
  AND2_X1 U473 ( .A1(n360), .A2(n455), .ZN(n702) );
  NAND2_X1 U474 ( .A1(n361), .A2(KEYINPUT44), .ZN(n597) );
  XNOR2_X1 U475 ( .A(n361), .B(G122), .ZN(n717) );
  XNOR2_X2 U476 ( .A(n399), .B(KEYINPUT35), .ZN(n361) );
  XNOR2_X1 U477 ( .A(n446), .B(n447), .ZN(n363) );
  NAND2_X1 U478 ( .A1(n574), .A2(n575), .ZN(n586) );
  NAND2_X1 U479 ( .A1(n562), .A2(n558), .ZN(n547) );
  NAND2_X1 U480 ( .A1(n574), .A2(n572), .ZN(n573) );
  NAND2_X1 U481 ( .A1(n364), .A2(n410), .ZN(n405) );
  NAND2_X1 U482 ( .A1(n409), .A2(n407), .ZN(n364) );
  NAND2_X1 U483 ( .A1(n404), .A2(n352), .ZN(n403) );
  AND2_X1 U484 ( .A1(n598), .A2(n599), .ZN(n600) );
  BUF_X1 U485 ( .A(n562), .Z(n366) );
  XNOR2_X2 U486 ( .A(n382), .B(n448), .ZN(n562) );
  NOR2_X2 U487 ( .A1(n681), .A2(n696), .ZN(n682) );
  XNOR2_X1 U488 ( .A(n367), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U489 ( .A1(n368), .A2(n418), .ZN(n378) );
  XNOR2_X1 U490 ( .A(n607), .B(n356), .ZN(n368) );
  NAND2_X1 U491 ( .A1(n576), .A2(n640), .ZN(n616) );
  XNOR2_X1 U492 ( .A(n370), .B(n369), .ZN(G75) );
  NAND2_X1 U493 ( .A1(n674), .A2(n427), .ZN(n370) );
  XNOR2_X1 U494 ( .A(n548), .B(KEYINPUT36), .ZN(n372) );
  INV_X1 U495 ( .A(n478), .ZN(n374) );
  NOR2_X1 U496 ( .A1(n549), .A2(n630), .ZN(n404) );
  XNOR2_X1 U497 ( .A(n378), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X2 U498 ( .A(n379), .B(n422), .ZN(n591) );
  NAND2_X1 U499 ( .A1(n381), .A2(n380), .ZN(n399) );
  INV_X1 U500 ( .A(n477), .ZN(n434) );
  XNOR2_X2 U501 ( .A(n446), .B(G134), .ZN(n513) );
  NAND2_X1 U502 ( .A1(n384), .A2(n383), .ZN(n637) );
  NAND2_X1 U503 ( .A1(n385), .A2(n392), .ZN(n383) );
  NOR2_X1 U504 ( .A1(n387), .A2(n386), .ZN(n384) );
  NAND2_X1 U505 ( .A1(n392), .A2(n389), .ZN(n542) );
  INV_X1 U506 ( .A(n467), .ZN(n391) );
  NAND2_X1 U507 ( .A1(n467), .A2(n396), .ZN(n395) );
  NAND2_X2 U508 ( .A1(n603), .A2(KEYINPUT2), .ZN(n633) );
  XNOR2_X2 U509 ( .A(n434), .B(n435), .ZN(n467) );
  NOR2_X1 U510 ( .A1(n400), .A2(n622), .ZN(n623) );
  NOR2_X1 U511 ( .A1(n400), .A2(n617), .ZN(n619) );
  NAND2_X1 U512 ( .A1(n405), .A2(n403), .ZN(n565) );
  NAND2_X1 U513 ( .A1(n408), .A2(n556), .ZN(n407) );
  INV_X1 U514 ( .A(n556), .ZN(n411) );
  INV_X1 U515 ( .A(n554), .ZN(n412) );
  XNOR2_X2 U516 ( .A(n413), .B(n465), .ZN(n640) );
  NAND2_X1 U517 ( .A1(n596), .A2(KEYINPUT44), .ZN(n415) );
  NOR2_X1 U518 ( .A1(n595), .A2(n608), .ZN(n416) );
  NOR2_X2 U519 ( .A1(n587), .A2(n640), .ZN(n608) );
  XNOR2_X1 U520 ( .A(n417), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U521 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U522 ( .A(n420), .B(n605), .ZN(n419) );
  XNOR2_X1 U523 ( .A(n686), .B(n685), .ZN(n687) );
  BUF_X1 U524 ( .A(n688), .Z(n692) );
  AND2_X1 U525 ( .A1(n349), .A2(n673), .ZN(n427) );
  AND2_X1 U526 ( .A1(n495), .A2(G210), .ZN(n428) );
  INV_X1 U527 ( .A(KEYINPUT105), .ZN(n577) );
  XNOR2_X1 U528 ( .A(n475), .B(n428), .ZN(n476) );
  INV_X1 U529 ( .A(G469), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n555), .B(KEYINPUT66), .ZN(n556) );
  XNOR2_X1 U531 ( .A(n479), .B(G472), .ZN(n480) );
  XNOR2_X1 U532 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U533 ( .A(n684), .B(n683), .ZN(n685) );
  INV_X1 U534 ( .A(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U535 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n437) );
  XNOR2_X1 U536 ( .A(G101), .B(G110), .ZN(n429) );
  XNOR2_X1 U537 ( .A(n350), .B(n429), .ZN(n444) );
  XOR2_X1 U538 ( .A(n454), .B(KEYINPUT90), .Z(n431) );
  NAND2_X1 U539 ( .A1(G227), .A2(n455), .ZN(n430) );
  XNOR2_X1 U540 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U541 ( .A(n444), .B(n432), .ZN(n435) );
  XOR2_X2 U542 ( .A(G143), .B(G128), .Z(n446) );
  XNOR2_X1 U543 ( .A(n467), .B(KEYINPUT57), .ZN(n436) );
  XNOR2_X1 U544 ( .A(n437), .B(n436), .ZN(n605) );
  XOR2_X1 U545 ( .A(KEYINPUT87), .B(KEYINPUT75), .Z(n439) );
  NAND2_X1 U546 ( .A1(G210), .A2(n471), .ZN(n438) );
  XNOR2_X1 U547 ( .A(n439), .B(n438), .ZN(n448) );
  NAND2_X1 U548 ( .A1(G224), .A2(n455), .ZN(n441) );
  XOR2_X1 U549 ( .A(n442), .B(n453), .Z(n447) );
  XNOR2_X1 U550 ( .A(n562), .B(KEYINPUT38), .ZN(n653) );
  INV_X1 U551 ( .A(n602), .ZN(n449) );
  NAND2_X1 U552 ( .A1(n449), .A2(G234), .ZN(n451) );
  XNOR2_X1 U553 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n450) );
  XNOR2_X1 U554 ( .A(n451), .B(n450), .ZN(n463) );
  NAND2_X1 U555 ( .A1(G221), .A2(n463), .ZN(n452) );
  XNOR2_X1 U556 ( .A(KEYINPUT21), .B(n452), .ZN(n639) );
  XNOR2_X1 U557 ( .A(n453), .B(KEYINPUT10), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n454), .B(n496), .ZN(n706) );
  NAND2_X1 U559 ( .A1(n455), .A2(G234), .ZN(n457) );
  XNOR2_X1 U560 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n456) );
  XNOR2_X1 U561 ( .A(n706), .B(n462), .ZN(n694) );
  NOR2_X1 U562 ( .A1(G902), .A2(n694), .ZN(n465) );
  NAND2_X1 U563 ( .A1(G217), .A2(n463), .ZN(n464) );
  XOR2_X1 U564 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n466) );
  XNOR2_X1 U565 ( .A(KEYINPUT94), .B(n470), .ZN(n592) );
  NAND2_X1 U566 ( .A1(G214), .A2(n471), .ZN(n472) );
  XOR2_X1 U567 ( .A(KEYINPUT88), .B(n472), .Z(n652) );
  XNOR2_X1 U568 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U569 ( .A1(G953), .A2(G237), .ZN(n495) );
  NOR2_X1 U570 ( .A1(n606), .A2(G902), .ZN(n481) );
  XNOR2_X1 U571 ( .A(KEYINPUT96), .B(KEYINPUT70), .ZN(n479) );
  NOR2_X1 U572 ( .A1(n652), .A2(n543), .ZN(n482) );
  XOR2_X1 U573 ( .A(KEYINPUT30), .B(n482), .Z(n483) );
  NAND2_X1 U574 ( .A1(G234), .A2(G237), .ZN(n484) );
  XNOR2_X1 U575 ( .A(n484), .B(KEYINPUT14), .ZN(n485) );
  NAND2_X1 U576 ( .A1(G952), .A2(n485), .ZN(n667) );
  NOR2_X1 U577 ( .A1(G953), .A2(n667), .ZN(n571) );
  NAND2_X1 U578 ( .A1(G902), .A2(n485), .ZN(n569) );
  OR2_X1 U579 ( .A1(n455), .A2(n569), .ZN(n486) );
  XNOR2_X1 U580 ( .A(KEYINPUT106), .B(n486), .ZN(n487) );
  NOR2_X1 U581 ( .A1(G900), .A2(n487), .ZN(n488) );
  NOR2_X1 U582 ( .A1(n571), .A2(n488), .ZN(n489) );
  XOR2_X1 U583 ( .A(KEYINPUT76), .B(n489), .Z(n527) );
  NAND2_X1 U584 ( .A1(n490), .A2(n527), .ZN(n552) );
  XNOR2_X1 U585 ( .A(n492), .B(n491), .ZN(n524) );
  XOR2_X1 U586 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n494) );
  XNOR2_X1 U587 ( .A(KEYINPUT13), .B(G475), .ZN(n493) );
  XNOR2_X1 U588 ( .A(n494), .B(n493), .ZN(n512) );
  NAND2_X1 U589 ( .A1(G214), .A2(n495), .ZN(n498) );
  INV_X1 U590 ( .A(n496), .ZN(n497) );
  XNOR2_X1 U591 ( .A(n498), .B(n497), .ZN(n510) );
  XOR2_X1 U592 ( .A(G122), .B(G104), .Z(n500) );
  XNOR2_X1 U593 ( .A(n500), .B(n499), .ZN(n504) );
  XOR2_X1 U594 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n502) );
  XNOR2_X1 U595 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n504), .B(n503), .ZN(n508) );
  XOR2_X1 U597 ( .A(KEYINPUT98), .B(KEYINPUT101), .Z(n506) );
  XNOR2_X1 U598 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n505) );
  XNOR2_X1 U599 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U600 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n510), .B(n509), .ZN(n684) );
  NOR2_X1 U602 ( .A1(G902), .A2(n684), .ZN(n511) );
  XOR2_X1 U603 ( .A(n512), .B(n511), .Z(n522) );
  INV_X1 U604 ( .A(n513), .ZN(n520) );
  NAND2_X1 U605 ( .A1(G217), .A2(n514), .ZN(n515) );
  XNOR2_X1 U606 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U607 ( .A(n520), .B(n519), .ZN(n690) );
  NOR2_X1 U608 ( .A1(G902), .A2(n690), .ZN(n521) );
  XOR2_X1 U609 ( .A(G478), .B(n521), .Z(n551) );
  NAND2_X1 U610 ( .A1(n522), .A2(n551), .ZN(n617) );
  INV_X1 U611 ( .A(n617), .ZN(n627) );
  AND2_X1 U612 ( .A1(n524), .A2(n627), .ZN(n630) );
  INV_X1 U613 ( .A(n522), .ZN(n550) );
  INV_X1 U614 ( .A(n551), .ZN(n523) );
  NAND2_X1 U615 ( .A1(n550), .A2(n523), .ZN(n622) );
  INV_X1 U616 ( .A(n622), .ZN(n625) );
  NAND2_X1 U617 ( .A1(n524), .A2(n625), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n525), .B(KEYINPUT40), .ZN(n723) );
  INV_X1 U619 ( .A(n543), .ZN(n643) );
  INV_X1 U620 ( .A(n639), .ZN(n526) );
  XNOR2_X1 U621 ( .A(KEYINPUT67), .B(n528), .ZN(n544) );
  AND2_X1 U622 ( .A1(n643), .A2(n544), .ZN(n529) );
  XNOR2_X1 U623 ( .A(n529), .B(KEYINPUT28), .ZN(n530) );
  NAND2_X1 U624 ( .A1(n530), .A2(n542), .ZN(n536) );
  XOR2_X1 U625 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n532) );
  NOR2_X1 U626 ( .A1(n652), .A2(n653), .ZN(n658) );
  NAND2_X1 U627 ( .A1(n658), .A2(n654), .ZN(n531) );
  XNOR2_X1 U628 ( .A(n532), .B(n531), .ZN(n670) );
  NOR2_X1 U629 ( .A1(n536), .A2(n670), .ZN(n533) );
  XOR2_X1 U630 ( .A(KEYINPUT42), .B(n533), .Z(n718) );
  NAND2_X1 U631 ( .A1(n723), .A2(n718), .ZN(n535) );
  XNOR2_X1 U632 ( .A(KEYINPUT46), .B(KEYINPUT81), .ZN(n534) );
  XNOR2_X1 U633 ( .A(n535), .B(n534), .ZN(n541) );
  INV_X1 U634 ( .A(n652), .ZN(n558) );
  NOR2_X1 U635 ( .A1(n625), .A2(n627), .ZN(n538) );
  XNOR2_X1 U636 ( .A(KEYINPUT104), .B(n538), .ZN(n656) );
  XNOR2_X1 U637 ( .A(n539), .B(KEYINPUT47), .ZN(n540) );
  NAND2_X1 U638 ( .A1(n541), .A2(n540), .ZN(n549) );
  INV_X1 U639 ( .A(n637), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT6), .B(n543), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n544), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT109), .ZN(n546) );
  NOR2_X1 U643 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U644 ( .A(KEYINPUT110), .B(n348), .ZN(n720) );
  NAND2_X1 U645 ( .A1(n551), .A2(n550), .ZN(n582) );
  NOR2_X1 U646 ( .A1(n552), .A2(n582), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n366), .A2(n553), .ZN(n621) );
  XNOR2_X1 U648 ( .A(n621), .B(KEYINPUT78), .ZN(n554) );
  INV_X1 U649 ( .A(KEYINPUT48), .ZN(n555) );
  NAND2_X1 U650 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U651 ( .A(n559), .B(KEYINPUT107), .ZN(n560) );
  NAND2_X1 U652 ( .A1(n560), .A2(n575), .ZN(n561) );
  XNOR2_X1 U653 ( .A(n561), .B(KEYINPUT43), .ZN(n564) );
  INV_X1 U654 ( .A(n366), .ZN(n563) );
  NAND2_X1 U655 ( .A1(n564), .A2(n563), .ZN(n631) );
  NAND2_X1 U656 ( .A1(n565), .A2(n631), .ZN(n713) );
  NOR2_X1 U657 ( .A1(n585), .A2(n575), .ZN(n566) );
  NAND2_X1 U658 ( .A1(n640), .A2(n566), .ZN(n567) );
  XNOR2_X1 U659 ( .A(n567), .B(KEYINPUT73), .ZN(n572) );
  NOR2_X1 U660 ( .A1(G898), .A2(n455), .ZN(n568) );
  XNOR2_X1 U661 ( .A(KEYINPUT89), .B(n568), .ZN(n698) );
  NOR2_X1 U662 ( .A1(n569), .A2(n698), .ZN(n570) );
  NOR2_X1 U663 ( .A1(n643), .A2(n586), .ZN(n576) );
  XNOR2_X1 U664 ( .A(KEYINPUT83), .B(n596), .ZN(n584) );
  INV_X1 U665 ( .A(n591), .ZN(n580) );
  XNOR2_X1 U666 ( .A(n588), .B(n577), .ZN(n578) );
  NAND2_X1 U667 ( .A1(n578), .A2(n585), .ZN(n579) );
  XNOR2_X2 U668 ( .A(n579), .B(KEYINPUT33), .ZN(n672) );
  OR2_X1 U669 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n643), .A2(n588), .ZN(n648) );
  NOR2_X1 U671 ( .A1(n591), .A2(n648), .ZN(n590) );
  XNOR2_X1 U672 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n589) );
  XNOR2_X1 U673 ( .A(n590), .B(n589), .ZN(n628) );
  OR2_X1 U674 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U675 ( .A1(n643), .A2(n593), .ZN(n612) );
  NOR2_X1 U676 ( .A1(n628), .A2(n612), .ZN(n594) );
  NOR2_X1 U677 ( .A1(n656), .A2(n594), .ZN(n595) );
  XNOR2_X1 U678 ( .A(n597), .B(KEYINPUT82), .ZN(n598) );
  NOR2_X2 U679 ( .A1(n603), .A2(KEYINPUT2), .ZN(n632) );
  NOR2_X4 U680 ( .A1(n604), .A2(n632), .ZN(n688) );
  NAND2_X1 U681 ( .A1(n688), .A2(G472), .ZN(n607) );
  XNOR2_X1 U682 ( .A(G101), .B(n608), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U684 ( .A1(n612), .A2(n625), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n610), .B(KEYINPUT112), .ZN(n611) );
  XNOR2_X1 U686 ( .A(G104), .B(n611), .ZN(G6) );
  XOR2_X1 U687 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n614) );
  NAND2_X1 U688 ( .A1(n612), .A2(n627), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U690 ( .A(G107), .B(n615), .ZN(G9) );
  XNOR2_X1 U691 ( .A(n616), .B(G110), .ZN(G12) );
  XNOR2_X1 U692 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n620) );
  XOR2_X1 U694 ( .A(G128), .B(n620), .Z(G30) );
  XNOR2_X1 U695 ( .A(G143), .B(n621), .ZN(G45) );
  XOR2_X1 U696 ( .A(KEYINPUT114), .B(n623), .Z(n624) );
  XNOR2_X1 U697 ( .A(G146), .B(n624), .ZN(G48) );
  NAND2_X1 U698 ( .A1(n628), .A2(n625), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n626), .B(G113), .ZN(G15) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n629), .B(G116), .ZN(G18) );
  XOR2_X1 U702 ( .A(G134), .B(n630), .Z(G36) );
  XNOR2_X1 U703 ( .A(G140), .B(n631), .ZN(G42) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT77), .ZN(n634) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n635), .B(KEYINPUT80), .ZN(n674) );
  OR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT50), .B(n638), .ZN(n646) );
  XOR2_X1 U709 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n642) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(n644) );
  NOR2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U715 ( .A(KEYINPUT51), .B(n649), .ZN(n650) );
  NOR2_X1 U716 ( .A1(n670), .A2(n650), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT116), .B(n651), .Z(n664) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n660) );
  INV_X1 U720 ( .A(n656), .ZN(n657) );
  NAND2_X1 U721 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U722 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U723 ( .A(KEYINPUT117), .B(n661), .Z(n662) );
  NAND2_X1 U724 ( .A1(n672), .A2(n662), .ZN(n663) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U726 ( .A(KEYINPUT52), .B(n665), .Z(n666) );
  NOR2_X1 U727 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U728 ( .A(n668), .B(KEYINPUT118), .ZN(n669) );
  INV_X1 U729 ( .A(n670), .ZN(n671) );
  NAND2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U731 ( .A(KEYINPUT55), .B(KEYINPUT84), .Z(n676) );
  XNOR2_X1 U732 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n675) );
  XNOR2_X1 U733 ( .A(n676), .B(n675), .ZN(n677) );
  XOR2_X1 U734 ( .A(n678), .B(n677), .Z(n680) );
  NAND2_X1 U735 ( .A1(n688), .A2(G210), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U737 ( .A(n682), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U738 ( .A1(n688), .A2(G475), .ZN(n686) );
  XOR2_X1 U739 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n683) );
  NAND2_X1 U740 ( .A1(G478), .A2(n692), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U742 ( .A1(n696), .A2(n691), .ZN(G63) );
  NAND2_X1 U743 ( .A1(G217), .A2(n692), .ZN(n693) );
  XNOR2_X1 U744 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U745 ( .A1(n696), .A2(n695), .ZN(G66) );
  XNOR2_X1 U746 ( .A(n697), .B(KEYINPUT122), .ZN(n699) );
  NAND2_X1 U747 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n700) );
  XNOR2_X1 U749 ( .A(KEYINPUT61), .B(n700), .ZN(n701) );
  AND2_X1 U750 ( .A1(n701), .A2(G898), .ZN(n703) );
  NOR2_X1 U751 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U752 ( .A(n705), .B(n704), .ZN(G69) );
  XOR2_X1 U753 ( .A(n706), .B(KEYINPUT123), .Z(n707) );
  XNOR2_X1 U754 ( .A(n708), .B(n707), .ZN(n712) );
  XNOR2_X1 U755 ( .A(G227), .B(n712), .ZN(n709) );
  NAND2_X1 U756 ( .A1(n709), .A2(G900), .ZN(n710) );
  NAND2_X1 U757 ( .A1(n710), .A2(G953), .ZN(n711) );
  XNOR2_X1 U758 ( .A(n711), .B(KEYINPUT124), .ZN(n716) );
  XNOR2_X1 U759 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U760 ( .A1(n714), .A2(n455), .ZN(n715) );
  NAND2_X1 U761 ( .A1(n716), .A2(n715), .ZN(G72) );
  XNOR2_X1 U762 ( .A(n717), .B(KEYINPUT125), .ZN(G24) );
  XNOR2_X1 U763 ( .A(G137), .B(n718), .ZN(n719) );
  XNOR2_X1 U764 ( .A(n719), .B(KEYINPUT126), .ZN(G39) );
  XNOR2_X1 U765 ( .A(G125), .B(KEYINPUT37), .ZN(n721) );
  XNOR2_X1 U766 ( .A(n721), .B(n720), .ZN(G27) );
  XNOR2_X1 U767 ( .A(G119), .B(n722), .ZN(G21) );
  XNOR2_X1 U768 ( .A(G131), .B(n723), .ZN(G33) );
endmodule

