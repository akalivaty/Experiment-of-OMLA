//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  AND3_X1   g042(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n461), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OAI221_X1 g050(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n466), .A2(new_n470), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(G124), .A2(new_n478), .B1(new_n479), .B2(G136), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND3_X1   g057(.A1(new_n463), .A2(new_n465), .A3(G138), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n488), .A3(KEYINPUT70), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n463), .A2(new_n465), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n470), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(new_n470), .ZN(new_n497));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n462), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n495), .A2(new_n496), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n496), .B1(new_n495), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n506), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(G88), .A2(new_n514), .B1(new_n516), .B2(G50), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(new_n511), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n514), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT73), .B(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n520), .B(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n513), .A2(new_n530), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n508), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n508), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(G81), .A2(new_n514), .B1(new_n516), .B2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n538), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT9), .B1(new_n515), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n506), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n513), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n553), .A2(new_n561), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n514), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n506), .A2(G61), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(KEYINPUT77), .B1(G73), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n506), .A2(new_n572), .A3(G61), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n508), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n513), .A2(new_n575), .B1(new_n515), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(G85), .A2(new_n514), .B1(new_n516), .B2(G47), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n508), .B2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n514), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT78), .B(G66), .Z(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n555), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n516), .B2(G54), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n583), .B1(new_n590), .B2(G868), .ZN(G284));
  OAI21_X1  g166(.A(new_n583), .B1(new_n590), .B2(G868), .ZN(G321));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G299), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(G168), .ZN(G297));
  OAI21_X1  g170(.A(new_n594), .B1(new_n593), .B2(G168), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n597), .B2(G860), .ZN(G148));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n590), .A2(new_n597), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n543), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n599), .A3(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n472), .A2(new_n460), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(G2100), .Z(new_n611));
  OAI221_X1 g186(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n478), .A2(G123), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n479), .A2(G135), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G2096), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n617), .ZN(G156));
  XOR2_X1   g193(.A(G1341), .B(G1348), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT82), .ZN(new_n620));
  XOR2_X1   g195(.A(G2451), .B(G2454), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT16), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n620), .B(new_n622), .Z(new_n623));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n623), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT83), .Z(G401));
  INV_X1    g210(.A(KEYINPUT18), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(G2100), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(new_n616), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(G227));
  XNOR2_X1  g223(.A(G1961), .B(G1966), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT20), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n650), .A2(new_n652), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n659), .A2(new_n655), .A3(new_n653), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n657), .B(new_n660), .C1(new_n655), .C2(new_n659), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1991), .B(G1996), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G229));
  NOR2_X1   g244(.A1(G6), .A2(G16), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n578), .B2(G16), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT32), .B(G1981), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(G166), .A2(G16), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G16), .B2(G22), .ZN(new_n675));
  INV_X1    g250(.A(G1971), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n675), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G23), .ZN(new_n680));
  INV_X1    g255(.A(G288), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT33), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n671), .A2(new_n672), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n678), .A2(KEYINPUT34), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT86), .B(G29), .Z(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G25), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n479), .A2(G131), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT87), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n478), .A2(G119), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n466), .A2(G107), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT88), .Z(new_n696));
  INV_X1    g271(.A(new_n688), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n689), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(KEYINPUT34), .B1(new_n678), .B2(new_n686), .ZN(new_n701));
  MUX2_X1   g276(.A(G24), .B(G290), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n698), .B2(new_n699), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n687), .A2(new_n700), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT36), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n697), .A2(G35), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n697), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G2090), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n679), .A2(G20), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT23), .Z(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G299), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1956), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT96), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G33), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT90), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT25), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n479), .A2(G139), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n466), .B1(new_n723), .B2(KEYINPUT91), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(KEYINPUT91), .B2(new_n723), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n718), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G2072), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n688), .A2(G26), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n478), .A2(G128), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n466), .A2(G116), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n479), .A2(KEYINPUT89), .A3(G140), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT89), .B1(new_n479), .B2(G140), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n731), .B1(new_n732), .B2(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n730), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2067), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n728), .B(new_n738), .C1(new_n709), .C2(G2090), .ZN(new_n739));
  NOR2_X1   g314(.A1(G4), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n590), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G1348), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n717), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n478), .A2(G129), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n479), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT26), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(G105), .B2(new_n460), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n745), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n744), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n742), .A2(new_n743), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n679), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n543), .B2(new_n679), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1341), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n753), .A2(new_n754), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n741), .B2(G1348), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n755), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G168), .A2(new_n679), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n679), .B2(G21), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n717), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n615), .B2(new_n688), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT95), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n763), .B2(new_n764), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT24), .B(G34), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n688), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT93), .Z(new_n775));
  INV_X1    g350(.A(G160), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n717), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n679), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n679), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n765), .A2(new_n772), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n739), .A2(new_n761), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n727), .A2(G2072), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT92), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n697), .A2(G27), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n697), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2078), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n716), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n706), .A2(new_n791), .ZN(G150));
  INV_X1    g367(.A(G150), .ZN(G311));
  AOI22_X1  g368(.A1(G93), .A2(new_n514), .B1(new_n516), .B2(G55), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(new_n508), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n543), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n543), .A2(new_n797), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT38), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n590), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n807), .A2(new_n808), .A3(G860), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n799), .A2(G860), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT37), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(new_n811), .ZN(G145));
  XNOR2_X1  g387(.A(new_n481), .B(new_n776), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n615), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n495), .A2(new_n502), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n736), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n752), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(new_n726), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n726), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI221_X1 g396(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G130), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n479), .A2(G142), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(new_n609), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n695), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n814), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(KEYINPUT98), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(G37), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n814), .ZN(new_n832));
  INV_X1    g407(.A(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(new_n819), .A3(new_n818), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n834), .B2(new_n830), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(KEYINPUT99), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n837), .B(new_n832), .C1(new_n834), .C2(new_n830), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n831), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g415(.A1(new_n799), .A2(G868), .ZN(new_n841));
  XOR2_X1   g416(.A(G303), .B(G290), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n578), .B(G288), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n842), .B(new_n843), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT101), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT42), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT102), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n590), .A2(G299), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n590), .A2(G299), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(KEYINPUT100), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n590), .A2(G299), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(KEYINPUT41), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(new_n854), .A3(new_n849), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n850), .A2(new_n852), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n803), .B(new_n600), .ZN(new_n860));
  MUX2_X1   g435(.A(new_n857), .B(new_n859), .S(new_n860), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n847), .B(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n846), .A2(KEYINPUT102), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n593), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n841), .B1(new_n862), .B2(new_n864), .ZN(G295));
  AOI21_X1  g440(.A(new_n841), .B1(new_n862), .B2(new_n864), .ZN(G331));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n867));
  XNOR2_X1  g442(.A(G168), .B(G301), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n803), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n803), .A2(new_n868), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n853), .A3(new_n855), .ZN(new_n873));
  INV_X1    g448(.A(new_n844), .ZN(new_n874));
  INV_X1    g449(.A(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n859), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n874), .B1(new_n873), .B2(new_n877), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n867), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n858), .B1(new_n876), .B2(new_n854), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n848), .A2(new_n849), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n872), .A2(KEYINPUT41), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n885), .A3(new_n844), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(new_n878), .A3(new_n879), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n882), .B1(new_n867), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT44), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n880), .B2(new_n881), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n886), .A2(new_n878), .A3(new_n867), .A4(new_n879), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n890), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n889), .B1(new_n895), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g471(.A(G1384), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n815), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(G160), .A2(G40), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n736), .B(G2067), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n752), .B(G1996), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT106), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n699), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n696), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n736), .A2(G2067), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n695), .B(new_n908), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n907), .B1(new_n902), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(G290), .A2(G1986), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT126), .Z(new_n916));
  OR2_X1    g491(.A1(new_n916), .A2(KEYINPUT48), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(KEYINPUT48), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n902), .B1(new_n903), .B2(new_n752), .ZN(new_n920));
  INV_X1    g495(.A(new_n902), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n921), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n902), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n911), .A2(new_n919), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n815), .A2(KEYINPUT71), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n495), .A2(new_n496), .A3(new_n502), .ZN(new_n931));
  AOI21_X1  g506(.A(G1384), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT107), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G2084), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n897), .B1(new_n503), .B2(new_n504), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT50), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n495), .B2(new_n502), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n901), .B1(new_n939), .B2(new_n933), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(new_n935), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n942));
  INV_X1    g517(.A(G40), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n471), .A2(new_n474), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n942), .B(new_n944), .C1(new_n939), .C2(KEYINPUT45), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n936), .B2(new_n899), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n900), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n764), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT121), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n941), .A2(new_n948), .A3(KEYINPUT121), .ZN(new_n951));
  INV_X1    g526(.A(G8), .ZN(new_n952));
  NOR2_X1   g527(.A1(G168), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT122), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n950), .A2(new_n956), .A3(new_n951), .A4(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n951), .ZN(new_n959));
  OAI21_X1  g534(.A(G168), .B1(new_n959), .B2(new_n949), .ZN(new_n960));
  AND2_X1   g535(.A1(KEYINPUT51), .A2(G8), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n941), .A2(new_n948), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G8), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n953), .A2(KEYINPUT51), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n960), .A2(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT62), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n934), .A2(new_n938), .A3(new_n940), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n782), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n936), .A2(new_n899), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n939), .A2(KEYINPUT45), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n944), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n972), .B2(G2078), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n969), .A2(G2078), .ZN(new_n975));
  OR3_X1    g550(.A1(new_n946), .A2(new_n947), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G301), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n676), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT108), .B(G2090), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n967), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(G8), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n939), .A2(new_n944), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n991), .B(new_n993), .C1(new_n992), .C2(G288), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n990), .B1(G1976), .B2(new_n681), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n578), .B(G1981), .Z(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT110), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G305), .A2(G1981), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT49), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n997), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n933), .B(new_n897), .C1(new_n503), .C2(new_n504), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n901), .B1(new_n898), .B2(KEYINPUT50), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n972), .A2(new_n676), .B1(new_n1012), .B2(new_n979), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n986), .B1(new_n1013), .B2(new_n952), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n988), .A2(new_n1008), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n966), .A2(new_n977), .A3(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n958), .A2(new_n965), .A3(KEYINPUT62), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT124), .ZN(new_n1020));
  AOI211_X1 g595(.A(G1976), .B(G288), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n991), .B1(new_n1021), .B2(new_n1001), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n981), .A2(G8), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n987), .A3(new_n1008), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1008), .B1(new_n1023), .B2(new_n987), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT112), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n1008), .C1(new_n1023), .C2(new_n987), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n963), .A2(G286), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT63), .A3(new_n988), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1015), .A2(G286), .A3(new_n963), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1035), .A2(KEYINPUT63), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1025), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n970), .A2(new_n944), .A3(new_n971), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1956), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1011), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n560), .A2(KEYINPUT113), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n552), .B1(new_n560), .B2(KEYINPUT113), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n553), .A2(KEYINPUT57), .A3(new_n561), .A4(new_n562), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n989), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n939), .A2(new_n944), .A3(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G2067), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n967), .A2(new_n743), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n590), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1050), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1039), .A2(new_n1041), .A3(new_n1048), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1039), .A2(new_n1041), .A3(KEYINPUT114), .A4(new_n1048), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1050), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1048), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT118), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT117), .B(KEYINPUT61), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1059), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1073), .A2(new_n1068), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n901), .A2(G1996), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n971), .B(new_n1076), .C1(new_n932), .C2(KEYINPUT45), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND3_X1  g654(.A1(new_n1052), .A2(new_n1053), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n543), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT59), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT116), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1081), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n543), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1075), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1072), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1056), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT120), .B(new_n590), .C1(new_n1056), .C2(KEYINPUT60), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n967), .A2(new_n743), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1057), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1094), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1056), .A2(KEYINPUT60), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1092), .A2(new_n1093), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1072), .A2(new_n1091), .A3(KEYINPUT119), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1065), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n471), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n471), .A2(new_n1106), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n474), .A2(new_n943), .A3(new_n975), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(new_n900), .A3(new_n971), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n968), .A2(new_n973), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n968), .A2(new_n973), .A3(new_n976), .A4(G301), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1114), .A2(KEYINPUT54), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1015), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1112), .A2(G171), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n977), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1116), .B(new_n1119), .C1(new_n958), .C2(new_n965), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1020), .B(new_n1037), .C1(new_n1105), .C2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1050), .A2(KEYINPUT61), .A3(new_n1059), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1089), .B1(new_n1088), .B2(new_n543), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n800), .C1(new_n1087), .C2(new_n1081), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1071), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT118), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1066), .B(new_n1048), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1129), .B2(new_n1063), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1093), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1104), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1120), .B1(new_n1133), .B2(new_n1064), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1032), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1035), .A2(KEYINPUT63), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1024), .B(new_n1022), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT124), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1019), .B1(new_n1121), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n1140));
  NAND2_X1  g715(.A1(G290), .A2(G1986), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(new_n921), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT105), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n913), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n929), .B1(new_n1139), .B2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g721(.A(G319), .ZN(new_n1148));
  NOR3_X1   g722(.A1(G401), .A2(new_n1148), .A3(G227), .ZN(new_n1149));
  OAI21_X1  g723(.A(new_n1149), .B1(new_n667), .B2(new_n668), .ZN(new_n1150));
  INV_X1    g724(.A(new_n1150), .ZN(new_n1151));
  AND2_X1   g725(.A1(new_n839), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g726(.A(new_n1152), .B(KEYINPUT127), .C1(new_n893), .C2(new_n894), .ZN(new_n1153));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n839), .A2(new_n1151), .ZN(new_n1155));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n895), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g730(.A1(new_n1153), .A2(new_n1156), .ZN(G308));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(G225));
endmodule


