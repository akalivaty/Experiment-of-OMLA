//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  OAI211_X1 g001(.A(KEYINPUT69), .B(G134gat), .C1(new_n202), .C2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n204), .B(new_n205), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n203), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n203), .B2(new_n210), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT79), .B(G155gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT80), .B(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G148gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT78), .B1(new_n218), .B2(G141gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(G148gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n219), .B(new_n222), .C1(new_n221), .C2(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n217), .B(new_n223), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(KEYINPUT77), .B2(new_n224), .ZN(new_n228));
  XNOR2_X1  g027(.A(G141gat), .B(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT77), .ZN(new_n231));
  OAI221_X1 g030(.A(new_n228), .B1(KEYINPUT77), .B2(new_n224), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT84), .B1(new_n235), .B2(KEYINPUT4), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n212), .A2(new_n213), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n214), .A2(new_n234), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT82), .B1(new_n237), .B2(new_n233), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n236), .B(new_n241), .C1(new_n245), .C2(new_n240), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n233), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n237), .A2(KEYINPUT81), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n212), .B2(new_n213), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n246), .A2(new_n247), .A3(new_n248), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n243), .A2(new_n240), .A3(new_n244), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n248), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n248), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n234), .B1(new_n251), .B2(new_n253), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n245), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(KEYINPUT5), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G1gat), .B(G29gat), .Z(new_n265));
  XNOR2_X1  g064(.A(G57gat), .B(G85gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n263), .A3(new_n269), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  INV_X1    g075(.A(G218gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(KEYINPUT22), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G211gat), .B(G218gat), .Z(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n279), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n283), .B(KEYINPUT72), .Z(new_n284));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n287), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n297), .B2(new_n293), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT65), .B(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n300), .B2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n296), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT25), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n302), .A2(KEYINPUT25), .B1(new_n292), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n309), .B(KEYINPUT68), .Z(new_n310));
  INV_X1    g109(.A(new_n306), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n291), .B1(KEYINPUT26), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n297), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n296), .B1(new_n295), .B2(KEYINPUT27), .ZN(new_n317));
  AOI211_X1 g116(.A(new_n316), .B(new_n317), .C1(KEYINPUT27), .C2(new_n295), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n299), .A2(KEYINPUT27), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n317), .B1(new_n319), .B2(KEYINPUT66), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n305), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n284), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT28), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n313), .B(new_n314), .C1(new_n327), .C2(new_n318), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n283), .B1(new_n328), .B2(new_n305), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n282), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT73), .ZN(new_n331));
  XOR2_X1   g130(.A(G8gat), .B(G36gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT74), .ZN(new_n333));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n282), .C1(new_n326), .C2(new_n329), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n324), .A2(new_n325), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n339), .A2(new_n283), .B1(new_n284), .B2(new_n324), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n279), .B(new_n280), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n331), .A2(new_n336), .A3(new_n338), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n274), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT37), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n346), .A3(new_n338), .A4(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n335), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n330), .A2(KEYINPUT73), .B1(new_n340), .B2(new_n341), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n349), .B2(new_n338), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT38), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT88), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT88), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n353), .B(KEYINPUT38), .C1(new_n348), .C2(new_n350), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n346), .B1(new_n340), .B2(new_n282), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n341), .B1(new_n326), .B2(new_n329), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT38), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n347), .A3(new_n335), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n345), .A2(new_n352), .A3(new_n354), .A4(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT31), .B(G50gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n325), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT3), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n282), .A2(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT86), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n234), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n325), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n282), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(G228gat), .B(G233gat), .C1(new_n367), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT85), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n249), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n362), .A2(KEYINPUT85), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n233), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n369), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n361), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(G22gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n371), .A2(new_n377), .A3(new_n361), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n381), .ZN(new_n384));
  INV_X1    g183(.A(new_n382), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT40), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n248), .B1(new_n246), .B2(new_n255), .ZN(new_n389));
  OR3_X1    g188(.A1(new_n245), .A2(new_n261), .A3(new_n260), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT39), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n269), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n388), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n246), .A2(new_n255), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n260), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(KEYINPUT39), .A3(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n394), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(KEYINPUT40), .A3(new_n269), .A4(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n396), .A2(new_n401), .A3(new_n271), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n343), .A2(new_n403), .A3(KEYINPUT30), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT30), .B1(new_n343), .B2(new_n403), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  AOI211_X1 g205(.A(new_n406), .B(new_n336), .C1(new_n349), .C2(new_n338), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n331), .A2(new_n338), .A3(new_n342), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT75), .B1(new_n408), .B2(new_n335), .ZN(new_n409));
  OAI22_X1  g208(.A1(new_n404), .A2(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n387), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n359), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT36), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n324), .A2(new_n214), .ZN(new_n417));
  INV_X1    g216(.A(G227gat), .ZN(new_n418));
  INV_X1    g217(.A(G233gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n328), .A2(new_n305), .A3(new_n237), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n422), .B2(KEYINPUT32), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n422), .A2(KEYINPUT70), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT70), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n422), .B(KEYINPUT32), .C1(new_n424), .C2(new_n416), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n420), .B1(new_n417), .B2(new_n421), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT34), .B(new_n420), .C1(new_n417), .C2(new_n421), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(new_n434), .A3(new_n428), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n413), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n428), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n422), .A2(KEYINPUT70), .A3(new_n424), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n444), .B2(new_n423), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT71), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n436), .A2(new_n437), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT71), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n438), .B1(new_n448), .B2(new_n413), .ZN(new_n449));
  INV_X1    g248(.A(new_n405), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n343), .A2(new_n403), .A3(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n408), .A2(new_n335), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n406), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n408), .A2(KEYINPUT75), .A3(new_n335), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n274), .A2(new_n344), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n387), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n412), .A2(new_n449), .A3(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n427), .A2(new_n434), .A3(new_n428), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n434), .B1(new_n427), .B2(new_n428), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n387), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT90), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n465));
  NOR4_X1   g264(.A1(new_n460), .A2(new_n387), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT35), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(KEYINPUT35), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n457), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n274), .A2(new_n344), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT89), .B1(new_n410), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n463), .A3(new_n448), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G155gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G183gat), .B(G211gat), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n479), .B(new_n480), .Z(new_n481));
  XOR2_X1   g280(.A(G57gat), .B(G64gat), .Z(new_n482));
  OR2_X1    g281(.A1(G71gat), .A2(G78gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT9), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n484), .B(new_n483), .C1(new_n489), .C2(new_n486), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT21), .ZN(new_n492));
  AND2_X1   g291(.A1(G231gat), .A2(G233gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G127gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(KEYINPUT101), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n488), .A2(new_n490), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT101), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT21), .ZN(new_n501));
  INV_X1    g300(.A(G1gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT16), .ZN(new_n503));
  INV_X1    g302(.A(G22gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G15gat), .ZN(new_n505));
  INV_X1    g304(.A(G15gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G22gat), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT96), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT96), .B1(new_n505), .B2(new_n507), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n506), .A2(G22gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n504), .A2(G15gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT96), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n502), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n512), .A2(new_n519), .A3(G8gat), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n510), .B(new_n518), .C1(new_n511), .C2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n501), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n495), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n495), .A2(new_n524), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n481), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  INV_X1    g328(.A(new_n481), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G190gat), .B(G218gat), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536));
  INV_X1    g335(.A(G50gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(G43gat), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G43gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(G29gat), .A2(G36gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(G29gat), .A3(G36gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n538), .A2(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n539), .A3(G50gat), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT91), .B1(new_n539), .B2(G50gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n537), .A2(G43gat), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n536), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NOR3_X1   g351(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556));
  INV_X1    g355(.A(G29gat), .ZN(new_n557));
  INV_X1    g356(.A(G36gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n535), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n552), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(KEYINPUT94), .A3(new_n550), .A4(new_n545), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n538), .A2(new_n540), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n552), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n541), .B1(new_n570), .B2(new_n553), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(KEYINPUT17), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT7), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n574), .B2(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n583), .A3(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n562), .A2(new_n566), .B1(new_n571), .B2(new_n569), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT95), .B(KEYINPUT17), .Z(new_n589));
  OAI211_X1 g388(.A(new_n573), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n572), .ZN(new_n591));
  INV_X1    g390(.A(new_n587), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n591), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n534), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n597));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n534), .A3(new_n594), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n586), .A2(KEYINPUT102), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n587), .A2(new_n491), .A3(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n586), .B(new_n585), .C1(new_n497), .C2(KEYINPUT102), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n586), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n496), .B2(new_n499), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n604), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n604), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n614), .A3(new_n609), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n532), .A2(new_n603), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n523), .B(new_n573), .C1(new_n588), .C2(new_n589), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n520), .A2(new_n522), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n591), .A2(new_n628), .A3(KEYINPUT98), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT98), .B1(new_n591), .B2(new_n628), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n626), .B(new_n627), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT99), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n523), .B2(new_n588), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n591), .A2(new_n628), .A3(KEYINPUT98), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n627), .A4(new_n626), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n636), .A2(KEYINPUT18), .A3(new_n627), .A4(new_n626), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n523), .A2(new_n588), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n629), .B2(new_n630), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n627), .B(KEYINPUT13), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G197gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT11), .B(G169gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n640), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n640), .B2(new_n646), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n625), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n477), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n472), .A2(KEYINPUT104), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n472), .A2(KEYINPUT104), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT105), .B(G1gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n657), .A2(new_n455), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT106), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(KEYINPUT106), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(G8gat), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n669), .B1(new_n666), .B2(new_n667), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n668), .B(new_n672), .C1(new_n673), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n657), .B2(new_n449), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n448), .A2(new_n506), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n657), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n657), .A2(new_n463), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT107), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n477), .A2(new_n682), .A3(new_n603), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n477), .A2(new_n682), .A3(KEYINPUT44), .A4(new_n603), .ZN(new_n686));
  INV_X1    g485(.A(new_n532), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(new_n654), .A3(new_n624), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n685), .A2(new_n660), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G29gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n661), .A2(G29gat), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n477), .A2(new_n603), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n690), .A2(KEYINPUT109), .A3(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1328gat));
  INV_X1    g497(.A(new_n603), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n467), .A2(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n459), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(new_n688), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n558), .A3(new_n410), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND4_X1   g504(.A1(new_n410), .A2(new_n685), .A3(new_n686), .A4(new_n688), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n558), .B2(new_n706), .ZN(G1329gat));
  INV_X1    g506(.A(new_n449), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n685), .A2(new_n708), .A3(new_n686), .A4(new_n688), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n539), .A2(KEYINPUT111), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  INV_X1    g511(.A(new_n448), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(KEYINPUT111), .A3(G43gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n702), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n711), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n711), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1330gat));
  NAND4_X1  g517(.A1(new_n685), .A2(new_n387), .A3(new_n686), .A4(new_n688), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G50gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n537), .A3(new_n387), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(KEYINPUT48), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1331gat));
  INV_X1    g525(.A(new_n624), .ZN(new_n727));
  NOR4_X1   g526(.A1(new_n655), .A2(new_n532), .A3(new_n603), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n477), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n660), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g531(.A1(new_n729), .A2(KEYINPUT112), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n477), .A2(new_n734), .A3(new_n728), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n736), .B(new_n410), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n736), .A2(new_n410), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n737), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n730), .B2(new_n448), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n729), .A2(KEYINPUT113), .A3(new_n713), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n733), .A2(new_n708), .A3(new_n735), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G71gat), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n747), .B1(new_n746), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n387), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g553(.A1(new_n655), .A2(new_n687), .A3(new_n727), .ZN(new_n755));
  AND4_X1   g554(.A1(new_n660), .A2(new_n685), .A3(new_n686), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n655), .A2(new_n687), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n701), .B2(new_n757), .ZN(new_n758));
  AND4_X1   g557(.A1(KEYINPUT51), .A2(new_n477), .A3(new_n603), .A4(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n660), .A2(new_n574), .A3(new_n624), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n756), .A2(new_n574), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  NAND4_X1  g561(.A1(new_n685), .A2(new_n410), .A3(new_n686), .A4(new_n755), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n455), .A2(G92gat), .A3(new_n727), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n758), .B2(new_n759), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT52), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n764), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1337gat));
  AND4_X1   g570(.A1(new_n708), .A2(new_n685), .A3(new_n686), .A4(new_n755), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT114), .B(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n448), .A2(new_n624), .A3(new_n773), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n772), .A2(new_n773), .B1(new_n760), .B2(new_n774), .ZN(G1338gat));
  NAND4_X1  g574(.A1(new_n685), .A2(new_n387), .A3(new_n686), .A4(new_n755), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n463), .A2(G106gat), .A3(new_n727), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n758), .B2(new_n759), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT115), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT53), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(G106gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n783), .A4(new_n779), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(G1339gat));
  AND2_X1   g584(.A1(new_n625), .A2(new_n654), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787));
  INV_X1    g586(.A(new_n627), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n591), .A2(new_n628), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n634), .B2(new_n635), .ZN(new_n791));
  INV_X1    g590(.A(new_n644), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n650), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n643), .A2(new_n644), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n627), .B1(new_n636), .B2(new_n626), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT117), .B(new_n650), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n640), .A2(new_n646), .A3(new_n651), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(new_n800), .A3(new_n624), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n802), .B(new_n604), .C1(new_n610), .C2(new_n612), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n613), .A2(KEYINPUT54), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n610), .A2(new_n604), .A3(new_n612), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n620), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n621), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n803), .A2(new_n620), .ZN(new_n809));
  INV_X1    g608(.A(new_n612), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n608), .A2(new_n609), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n810), .B(new_n614), .C1(new_n811), .C2(new_n606), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(KEYINPUT54), .A3(new_n613), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT55), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n808), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n651), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n632), .A2(new_n638), .A3(new_n639), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n641), .A2(new_n645), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n818), .B1(new_n822), .B2(new_n800), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n699), .B1(new_n801), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n808), .A2(new_n816), .A3(new_n817), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n603), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n799), .A2(new_n800), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n786), .B1(new_n830), .B2(new_n532), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n661), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n464), .A2(new_n466), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n410), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n655), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n660), .A2(new_n455), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n448), .A2(new_n463), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n831), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n654), .A2(new_n206), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(G1340gat));
  INV_X1    g641(.A(new_n840), .ZN(new_n843));
  OAI21_X1  g642(.A(G120gat), .B1(new_n843), .B2(new_n727), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n624), .A2(new_n208), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT118), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n835), .B2(new_n846), .ZN(G1341gat));
  XOR2_X1   g646(.A(KEYINPUT69), .B(G127gat), .Z(new_n848));
  NOR3_X1   g647(.A1(new_n843), .A2(new_n532), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n836), .A2(new_n687), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT119), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n848), .ZN(G1342gat));
  NOR3_X1   g651(.A1(new_n835), .A2(G134gat), .A3(new_n699), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n843), .B2(new_n699), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NOR2_X1   g657(.A1(new_n838), .A2(new_n708), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n824), .A2(KEYINPUT120), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n825), .B1(new_n652), .B2(new_n653), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n799), .A2(new_n800), .A3(new_n624), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n603), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n829), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n532), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n625), .A2(new_n654), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n860), .B(new_n463), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n532), .B1(new_n864), .B2(new_n828), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n463), .B1(new_n870), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n859), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n655), .A2(G141gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n449), .A2(new_n387), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n831), .A2(new_n875), .A3(new_n661), .A4(new_n410), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(new_n655), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n873), .A2(new_n874), .B1(new_n877), .B2(G141gat), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n880), .B(G148gat), .C1(new_n873), .C2(new_n727), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT121), .B(new_n860), .C1(new_n831), .C2(new_n463), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n871), .B2(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n868), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .A3(new_n387), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n624), .A3(new_n859), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G148gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n882), .B1(new_n890), .B2(KEYINPUT59), .ZN(new_n891));
  AOI211_X1 g690(.A(KEYINPUT122), .B(new_n880), .C1(new_n889), .C2(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n881), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n218), .A3(new_n624), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1345gat));
  INV_X1    g694(.A(new_n215), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n873), .B2(new_n532), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n215), .A3(new_n687), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  NAND3_X1  g698(.A1(new_n876), .A2(new_n216), .A3(new_n603), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT123), .ZN(new_n901));
  INV_X1    g700(.A(new_n216), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n873), .B2(new_n699), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n660), .A2(new_n455), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT126), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(new_n463), .A3(new_n448), .A4(new_n886), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(new_n289), .A3(new_n654), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n831), .A2(new_n660), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT124), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n833), .A2(new_n455), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT125), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n655), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n908), .B1(new_n913), .B2(new_n289), .ZN(G1348gat));
  OAI21_X1  g713(.A(G176gat), .B1(new_n907), .B2(new_n727), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n624), .A2(new_n290), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n915), .B(KEYINPUT127), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(new_n300), .B1(new_n907), .B2(new_n532), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n295), .A2(KEYINPUT27), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n295), .A2(KEYINPUT27), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n687), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n916), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n923), .B(new_n929), .C1(new_n916), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  OR2_X1    g730(.A1(new_n907), .A2(new_n699), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(G190gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n932), .B2(G190gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n603), .A2(new_n296), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n934), .A2(new_n935), .B1(new_n916), .B2(new_n936), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n875), .A2(new_n455), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n910), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n655), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n906), .A2(new_n449), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(new_n888), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n655), .A2(G197gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n624), .A2(new_n946), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n939), .A2(KEYINPUT62), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT62), .B1(new_n939), .B2(new_n947), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n942), .A2(new_n624), .A3(new_n888), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n948), .B(new_n949), .C1(new_n946), .C2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n940), .A2(new_n276), .A3(new_n687), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n942), .A2(new_n687), .A3(new_n888), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n277), .A3(new_n603), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n943), .A2(new_n603), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n277), .ZN(G1355gat));
endmodule


