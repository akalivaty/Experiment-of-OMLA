//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT64), .A2(G137), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT11), .A2(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT66), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n194), .A2(new_n202), .A3(new_n197), .A4(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(G131), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G131), .B1(new_n198), .B2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n194), .A2(new_n197), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n194), .A2(new_n208), .A3(new_n197), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT71), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n204), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT0), .A3(G128), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n212), .A2(new_n214), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT64), .A2(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT64), .A2(G137), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n198), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n228), .B2(new_n195), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT11), .B1(new_n190), .B2(G134), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(new_n227), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n193), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n208), .B1(new_n233), .B2(new_n205), .ZN(new_n234));
  INV_X1    g048(.A(new_n209), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT72), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(new_n207), .B2(new_n209), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n217), .B2(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n216), .A2(new_n243), .A3(KEYINPUT1), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(G128), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n216), .A2(new_n218), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n246), .A2(KEYINPUT1), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n240), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n224), .A2(KEYINPUT30), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  INV_X1    g068(.A(G119), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n256), .A2(new_n258), .A3(G116), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n255), .B2(G116), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G119), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n254), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n254), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n258), .A3(G116), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n263), .A4(new_n260), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(KEYINPUT70), .B(new_n254), .C1(new_n259), .C2(new_n264), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n211), .A2(new_n223), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n238), .A2(new_n251), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n253), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  OR2_X1    g093(.A1(KEYINPUT73), .A2(G237), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT73), .A2(G237), .ZN(new_n281));
  AOI21_X1  g095(.A(G953), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G210), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT27), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G101), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g100(.A(new_n272), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n249), .B1(new_n246), .B2(new_n245), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n236), .B2(KEYINPUT72), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n289), .B2(new_n240), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(new_n224), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n278), .A2(new_n279), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n224), .A2(new_n272), .A3(new_n252), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n275), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n251), .A2(new_n210), .A3(new_n230), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n222), .B1(new_n204), .B2(new_n210), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n287), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT28), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n204), .A2(new_n213), .A3(new_n210), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n213), .B1(new_n204), .B2(new_n210), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(new_n222), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n251), .B1(new_n238), .B2(new_n239), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT72), .B(new_n229), .C1(new_n207), .C2(new_n209), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n272), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n302), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT76), .B(new_n302), .C1(new_n305), .C2(new_n308), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n301), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n292), .B1(new_n313), .B2(new_n286), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n278), .A2(new_n291), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT74), .B1(new_n315), .B2(KEYINPUT31), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n317), .B(new_n279), .C1(new_n278), .C2(new_n291), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n188), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n278), .A2(new_n293), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n284), .B(new_n285), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n324));
  AOI21_X1  g138(.A(G902), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n301), .A2(new_n324), .A3(new_n311), .A4(new_n312), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n322), .ZN(new_n327));
  INV_X1    g141(.A(new_n312), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT76), .B1(new_n293), .B2(new_n302), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n224), .A2(new_n252), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n293), .B1(new_n331), .B2(new_n272), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT28), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n324), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n325), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n320), .A2(KEYINPUT32), .B1(new_n335), .B2(G472), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n311), .A2(new_n312), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n290), .A2(new_n224), .B1(new_n297), .B2(new_n298), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n302), .B1(new_n339), .B2(new_n294), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n286), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n322), .B1(new_n305), .B2(new_n308), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n253), .B2(new_n277), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n317), .B1(new_n343), .B2(new_n279), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n279), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n315), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n341), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n187), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT77), .B(KEYINPUT32), .Z(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n337), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(KEYINPUT78), .B(new_n349), .C1(new_n347), .C2(new_n187), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n336), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  OR3_X1    g169(.A1(new_n355), .A2(KEYINPUT82), .A3(KEYINPUT16), .ZN(new_n356));
  XNOR2_X1  g170(.A(G125), .B(G140), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT82), .B1(new_n357), .B2(KEYINPUT16), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n355), .A2(KEYINPUT16), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n215), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n362));
  OAI211_X1 g176(.A(G146), .B(new_n356), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(KEYINPUT83), .A3(new_n215), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n256), .A2(new_n258), .A3(G128), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n255), .B2(G128), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT24), .B(G110), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n374));
  AOI21_X1  g188(.A(G128), .B1(new_n256), .B2(new_n258), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n373), .B2(KEYINPUT81), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G110), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n370), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n366), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n355), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT84), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n357), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n386), .A3(new_n215), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n363), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n377), .A2(new_n378), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n368), .A2(new_n369), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT22), .B(G137), .ZN(new_n393));
  INV_X1    g207(.A(G221), .ZN(new_n394));
  INV_X1    g208(.A(G234), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n395), .A3(G953), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n393), .B(new_n396), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n380), .A2(new_n392), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n397), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n366), .A2(new_n379), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  INV_X1    g215(.A(G902), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT25), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G217), .B1(new_n395), .B2(G902), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n398), .A2(KEYINPUT86), .A3(new_n401), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT86), .B1(new_n398), .B2(new_n401), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n395), .B2(G217), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G469), .ZN(new_n417));
  INV_X1    g231(.A(G953), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G227), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT87), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G140), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G104), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT3), .B1(new_n424), .B2(G107), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT3), .ZN(new_n426));
  INV_X1    g240(.A(G107), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(G104), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(G107), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(G101), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(G101), .ZN(new_n433));
  INV_X1    g247(.A(G101), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n425), .A2(new_n428), .A3(new_n434), .A4(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(KEYINPUT4), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n223), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n427), .A3(G104), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT88), .B1(new_n424), .B2(G107), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n427), .A2(G104), .ZN(new_n441));
  OAI211_X1 g255(.A(G101), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(new_n435), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n219), .B1(G128), .B2(new_n241), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n249), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT89), .B(KEYINPUT10), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n435), .A3(KEYINPUT10), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n251), .B2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n288), .A2(KEYINPUT90), .A3(new_n449), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n437), .B(new_n447), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n303), .A2(new_n304), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n423), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n442), .A2(new_n435), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n247), .A2(new_n250), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n445), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n458), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n212), .A2(new_n214), .A3(new_n458), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n437), .A2(new_n447), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT90), .B1(new_n288), .B2(new_n449), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n251), .A2(new_n448), .A3(new_n450), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n464), .B(new_n467), .C1(new_n304), .C2(new_n303), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n453), .A2(new_n454), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n423), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n417), .B(new_n402), .C1(new_n463), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(G469), .A2(G902), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n453), .A2(new_n454), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n422), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n469), .A3(new_n423), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n471), .B(new_n472), .C1(new_n417), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT9), .B(G234), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n394), .B1(new_n479), .B2(new_n402), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G214), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n270), .A2(new_n271), .A3(new_n432), .A4(new_n436), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n267), .A2(KEYINPUT5), .A3(new_n263), .A4(new_n260), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(G113), .C1(KEYINPUT5), .C2(new_n267), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n268), .A3(new_n443), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G122), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n495), .A3(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n288), .A2(new_n381), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n222), .A2(G125), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n418), .A2(G224), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n494), .A2(KEYINPUT91), .A3(new_n501), .A4(new_n496), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n288), .A2(KEYINPUT94), .A3(new_n381), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n222), .B2(G125), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n510), .A2(new_n513), .B1(new_n499), .B2(new_n512), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n490), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n443), .A2(new_n268), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n486), .A2(KEYINPUT93), .ZN(new_n518));
  OAI21_X1  g332(.A(G113), .B1(new_n267), .B2(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(KEYINPUT93), .B2(new_n486), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n443), .B1(new_n487), .B2(new_n268), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n493), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n402), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n506), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G210), .B1(G237), .B2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n506), .A2(new_n528), .A3(new_n526), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n484), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n482), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n280), .A2(new_n281), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(G214), .A3(new_n418), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT95), .B(G143), .Z(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n217), .A2(KEYINPUT95), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n282), .A2(G214), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n225), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT18), .A2(G131), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n357), .B(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n387), .B1(new_n545), .B2(new_n215), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n384), .A2(new_n386), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n215), .C1(new_n545), .C2(new_n548), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n537), .A2(new_n539), .A3(new_n225), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n550), .B(new_n363), .C1(new_n551), .C2(new_n540), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n424), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n547), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(G475), .A2(G902), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n559), .B(new_n225), .C1(new_n537), .C2(new_n539), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n551), .A2(new_n540), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n559), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n562), .B2(new_n366), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n556), .B(new_n557), .C1(new_n563), .C2(new_n555), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT20), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n547), .A2(new_n552), .A3(new_n555), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n364), .A2(new_n365), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n537), .A2(new_n539), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G131), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n537), .A2(new_n539), .A3(new_n225), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n559), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n560), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n547), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n574), .B2(new_n554), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT20), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n557), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n555), .A2(KEYINPUT97), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n563), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n578), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n402), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n565), .A2(new_n577), .B1(new_n582), .B2(G475), .ZN(new_n583));
  NAND2_X1  g397(.A1(G234), .A2(G237), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(G952), .A3(new_n418), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT21), .B(G898), .Z(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(G902), .A3(G953), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n248), .B2(G143), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n248), .A2(G143), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n217), .A2(G128), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n589), .ZN(new_n594));
  OAI21_X1  g408(.A(G134), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(G116), .B(G122), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n596), .A2(G107), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(G107), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n593), .A2(new_n591), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n198), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n595), .A2(new_n597), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT98), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n599), .A2(new_n198), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n600), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(KEYINPUT99), .A3(new_n600), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n262), .A2(G122), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n427), .B1(new_n608), .B2(KEYINPUT14), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n596), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n479), .A2(G217), .A3(new_n418), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n602), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G478), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n618), .A2(KEYINPUT15), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n402), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n619), .B1(new_n617), .B2(new_n402), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n583), .A2(new_n588), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n533), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n353), .A2(new_n416), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AND2_X1   g441(.A1(new_n416), .A2(new_n482), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n347), .B2(new_n402), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n320), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n602), .A2(new_n611), .A3(new_n615), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n615), .B1(new_n602), .B2(new_n611), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT33), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n614), .A2(new_n637), .A3(new_n616), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n638), .A3(G478), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n617), .A2(new_n618), .A3(new_n402), .ZN(new_n640));
  NAND2_X1  g454(.A1(G478), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n565), .A2(new_n577), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n402), .B1(new_n574), .B2(new_n578), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n563), .A2(new_n579), .ZN(new_n645));
  OAI21_X1  g459(.A(G475), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n642), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n532), .A2(KEYINPUT100), .A3(new_n588), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n528), .B1(new_n506), .B2(new_n526), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n529), .B(new_n525), .C1(new_n504), .C2(new_n505), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n483), .B(new_n588), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n647), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n633), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(new_n623), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n583), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n633), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n380), .A2(new_n392), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n399), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n413), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n409), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n314), .B2(new_n319), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n671), .B(new_n348), .C1(new_n672), .C2(new_n629), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n630), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .A3(new_n348), .A4(new_n671), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n677), .A3(new_n625), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT104), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT37), .B(G110), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  NAND3_X1  g495(.A1(new_n482), .A2(new_n532), .A3(new_n671), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n585), .B1(new_n587), .B2(G900), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n583), .A2(new_n661), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n353), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  NAND2_X1  g501(.A1(new_n530), .A2(new_n531), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT38), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n406), .A2(new_n408), .B1(new_n413), .B2(new_n669), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n483), .B1(new_n621), .B2(new_n622), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n583), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n684), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n482), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n693), .B1(KEYINPUT40), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n332), .A2(new_n322), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(G902), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n321), .A2(new_n322), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n629), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n320), .B2(KEYINPUT32), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n351), .B2(new_n352), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n696), .B(new_n702), .C1(KEYINPUT40), .C2(new_n695), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  AOI21_X1  g518(.A(KEYINPUT105), .B1(new_n647), .B2(new_n684), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n576), .B1(new_n575), .B2(new_n557), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n366), .A2(new_n571), .A3(new_n572), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n555), .B1(new_n707), .B2(new_n547), .ZN(new_n708));
  INV_X1    g522(.A(new_n557), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n708), .A2(KEYINPUT20), .A3(new_n566), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n646), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n642), .ZN(new_n712));
  AND4_X1   g526(.A1(KEYINPUT105), .A2(new_n711), .A3(new_n712), .A4(new_n684), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n353), .A2(new_n683), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT106), .B(G146), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G48));
  OAI21_X1  g531(.A(new_n402), .B1(new_n463), .B2(new_n470), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n471), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(KEYINPUT107), .A3(G469), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n480), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n655), .A2(new_n353), .A3(new_n416), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n353), .A2(new_n416), .A3(new_n663), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR2_X1   g542(.A1(new_n690), .A2(new_n624), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n532), .A3(new_n723), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n353), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  INV_X1    g546(.A(new_n723), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n688), .A2(new_n588), .A3(new_n692), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n330), .A2(new_n333), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n286), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n315), .B(new_n279), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n188), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n630), .A2(new_n415), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NAND2_X1  g556(.A1(new_n737), .A2(new_n738), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n187), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(new_n671), .C1(new_n629), .C2(new_n672), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n723), .A2(new_n532), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n711), .A2(new_n712), .A3(new_n684), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n647), .A2(KEYINPUT105), .A3(new_n684), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n745), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n381), .ZN(G27));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n335), .A2(G472), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n416), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n688), .A2(new_n484), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n482), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n754), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n650), .A2(new_n651), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n482), .A2(new_n483), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n751), .A3(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n336), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(KEYINPUT109), .A3(new_n416), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n764), .A2(new_n751), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n353), .A2(new_n771), .A3(new_n772), .A4(new_n416), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n765), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT78), .B1(new_n320), .B2(new_n349), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n348), .A2(new_n337), .A3(new_n350), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n415), .B1(new_n777), .B2(new_n336), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n771), .B1(new_n778), .B2(new_n772), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n770), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT110), .B(G131), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G33));
  INV_X1    g596(.A(new_n764), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n685), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  INV_X1    g599(.A(new_n760), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n583), .A2(new_n712), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT43), .Z(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(new_n671), .C1(new_n320), .C2(new_n630), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n476), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n474), .A2(KEYINPUT45), .A3(new_n475), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(G469), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n472), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n472), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT111), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(KEYINPUT111), .ZN(new_n800));
  OAI221_X1 g614(.A(new_n471), .B1(KEYINPUT46), .B2(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n481), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n694), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(new_n190), .ZN(G39));
  XOR2_X1   g619(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n802), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n714), .A2(new_n415), .A3(new_n760), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n353), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n354), .ZN(G42));
  NAND2_X1  g624(.A1(new_n721), .A2(new_n722), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n480), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n585), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n740), .A2(new_n788), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n760), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n723), .A2(new_n484), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT118), .Z(new_n818));
  INV_X1    g632(.A(new_n689), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n819), .A3(new_n815), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT50), .Z(new_n821));
  INV_X1    g635(.A(new_n702), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n786), .A2(new_n733), .A3(new_n585), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n416), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n711), .A3(new_n712), .ZN(new_n825));
  INV_X1    g639(.A(new_n745), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n823), .A2(new_n788), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n816), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(new_n416), .A3(new_n768), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  NAND2_X1  g648(.A1(new_n418), .A2(G952), .ZN(new_n835));
  INV_X1    g649(.A(new_n746), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n815), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n824), .B2(new_n653), .ZN(new_n838));
  OR4_X1    g652(.A1(new_n831), .A2(new_n832), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n653), .A2(new_n662), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n652), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n628), .A3(new_n631), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n626), .A2(new_n678), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n353), .A2(new_n416), .A3(new_n685), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n826), .A2(new_n714), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n623), .A2(new_n671), .A3(new_n583), .A4(new_n684), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n353), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n844), .B1(new_n783), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n353), .A2(new_n730), .B1(new_n740), .B2(new_n735), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n724), .A2(new_n851), .A3(new_n727), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n854), .A3(new_n780), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n682), .B1(new_n777), .B2(new_n336), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n752), .B1(new_n856), .B2(new_n685), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n661), .A2(new_n711), .A3(new_n483), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n763), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n482), .A2(new_n690), .A3(new_n684), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n702), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n715), .A4(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT115), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n826), .A2(new_n836), .A3(new_n714), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n686), .A2(new_n715), .A3(new_n861), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(KEYINPUT116), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n855), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n852), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n724), .A2(new_n851), .A3(new_n727), .A4(KEYINPUT113), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n850), .A2(new_n780), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n867), .A2(new_n862), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n853), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n880), .B(new_n853), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n872), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n850), .A2(new_n780), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n874), .A2(new_n875), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n867), .A2(new_n862), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n876), .B(KEYINPUT114), .Z(new_n890));
  XOR2_X1   g704(.A(new_n862), .B(KEYINPUT115), .Z(new_n891));
  INV_X1    g705(.A(new_n871), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n853), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n889), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n884), .B1(new_n894), .B2(new_n883), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n839), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n811), .B(KEYINPUT49), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n415), .A2(new_n484), .A3(new_n480), .A4(new_n787), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n819), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n702), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n418), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n882), .A2(new_n402), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(G210), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n494), .A2(new_n496), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n501), .ZN(new_n908));
  XOR2_X1   g722(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n902), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n904), .B2(new_n905), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n917), .B2(new_n910), .ZN(G51));
  INV_X1    g732(.A(new_n872), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n880), .B1(new_n888), .B2(new_n853), .ZN(new_n920));
  INV_X1    g734(.A(new_n881), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n884), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n472), .B(KEYINPUT57), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n470), .B2(new_n463), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n904), .A2(new_n796), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n901), .B1(new_n927), .B2(new_n928), .ZN(G54));
  INV_X1    g743(.A(KEYINPUT58), .ZN(new_n930));
  INV_X1    g744(.A(G475), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT121), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT121), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n903), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n575), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n901), .ZN(G60));
  AND2_X1   g752(.A1(new_n636), .A2(new_n638), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n641), .B(KEYINPUT59), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n924), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n895), .B2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n901), .ZN(G63));
  XNOR2_X1  g758(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT60), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n922), .A2(KEYINPUT122), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n882), .B2(new_n948), .ZN(new_n952));
  INV_X1    g766(.A(new_n412), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n902), .ZN(new_n955));
  INV_X1    g769(.A(new_n669), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n950), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n946), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n950), .A2(new_n952), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n669), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n902), .A3(new_n954), .A4(new_n945), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(G66));
  AOI21_X1  g776(.A(new_n418), .B1(new_n586), .B2(G224), .ZN(new_n963));
  INV_X1    g777(.A(new_n844), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n886), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n965), .B2(new_n418), .ZN(new_n966));
  INV_X1    g780(.A(G898), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n907), .B1(new_n967), .B2(G953), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G69));
  NAND2_X1  g783(.A1(G227), .A2(G900), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n780), .A2(new_n784), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n803), .A2(new_n763), .A3(new_n858), .A4(new_n759), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n809), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n804), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n857), .A2(new_n715), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n975), .A2(KEYINPUT125), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT125), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n972), .B(new_n974), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n418), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n418), .A2(G900), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n275), .A2(new_n276), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n253), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n549), .B1(new_n545), .B2(new_n548), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(G953), .B(new_n970), .C1(new_n985), .C2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n984), .A2(KEYINPUT127), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n981), .B2(new_n983), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n970), .A2(G953), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n786), .A2(new_n841), .A3(new_n695), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n804), .B1(new_n778), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n977), .A2(new_n703), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT62), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n999), .A2(new_n809), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n990), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n995), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n991), .A2(new_n1004), .ZN(G72));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT63), .ZN(new_n1007));
  INV_X1    g821(.A(new_n323), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n699), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n894), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n902), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1002), .A2(new_n322), .A3(new_n321), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n1008), .B2(new_n980), .ZN(new_n1014));
  INV_X1    g828(.A(new_n965), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n1010), .B(new_n1012), .C1(new_n1014), .C2(new_n1015), .ZN(G57));
endmodule


