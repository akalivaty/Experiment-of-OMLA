//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n468), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n468), .A2(new_n475), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G102), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(KEYINPUT70), .B2(KEYINPUT4), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n488), .B1(new_n493), .B2(new_n468), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n475), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n468), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n475), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n498), .A2(G2105), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT73), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n506), .B2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n503), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n504), .A2(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT71), .B(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(new_n507), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n509), .A2(new_n510), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT71), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT71), .A2(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT6), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n516), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n520), .A2(new_n521), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n518), .A2(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n514), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n532), .B1(new_n514), .B2(new_n528), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  AND2_X1   g111(.A1(new_n517), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  INV_X1    g113(.A(new_n526), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n513), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT75), .B(G90), .Z(new_n549));
  OAI22_X1  g124(.A1(new_n518), .A2(new_n548), .B1(new_n526), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n513), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n518), .A2(new_n554), .B1(new_n526), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n526), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT76), .B1(new_n511), .B2(new_n517), .ZN(new_n566));
  OAI21_X1  g141(.A(G91), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n517), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n525), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n520), .A2(new_n521), .A3(G65), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT77), .B1(new_n576), .B2(G651), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  AOI211_X1 g153(.A(new_n578), .B(new_n515), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT78), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n526), .A2(new_n564), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n511), .A2(new_n517), .A3(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G91), .B1(new_n571), .B2(new_n569), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n578), .B1(new_n586), .B2(new_n515), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n576), .A2(KEYINPUT77), .A3(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n581), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  NOR2_X1   g168(.A1(new_n565), .A2(new_n566), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT79), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n511), .A2(G74), .ZN(new_n597));
  AOI22_X1  g172(.A1(G651), .A2(new_n597), .B1(new_n537), .B2(G49), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n584), .A2(new_n599), .A3(G87), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(G288));
  NAND2_X1  g176(.A1(new_n584), .A2(G86), .ZN(new_n602));
  INV_X1    g177(.A(new_n513), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n520), .A2(new_n521), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n603), .A2(new_n607), .B1(new_n537), .B2(G48), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n602), .A2(new_n608), .ZN(G305));
  AOI22_X1  g184(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n513), .ZN(new_n611));
  INV_X1    g186(.A(G47), .ZN(new_n612));
  INV_X1    g187(.A(G85), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n518), .A2(new_n612), .B1(new_n526), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n611), .A2(new_n614), .ZN(G290));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  OR3_X1    g191(.A1(G171), .A2(KEYINPUT80), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT80), .B1(G171), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g193(.A(G92), .B1(new_n565), .B2(new_n566), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n605), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(G651), .A2(new_n623), .B1(new_n537), .B2(G54), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n584), .A2(new_n625), .A3(G92), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n617), .B(new_n618), .C1(new_n628), .C2(G868), .ZN(G284));
  XNOR2_X1  g204(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g205(.A1(G286), .A2(G868), .ZN(new_n631));
  XNOR2_X1  g206(.A(G299), .B(KEYINPUT82), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G297));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n628), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n645), .B(new_n647), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n484), .A2(G123), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n482), .A2(G135), .ZN(new_n650));
  NOR2_X1   g225(.A1(G99), .A2(G2105), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n653), .A2(G2096), .B1(new_n642), .B2(new_n643), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n648), .B(new_n654), .C1(G2096), .C2(new_n653), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2435), .ZN(new_n657));
  XOR2_X1   g232(.A(G2427), .B(G2438), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT14), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1341), .B(G1348), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2443), .B(G2446), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G14), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XOR2_X1   g246(.A(G2067), .B(G2678), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n671), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  AOI21_X1  g255(.A(KEYINPUT18), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n678), .B(new_n681), .Z(G227));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n693), .B(new_n694), .C1(new_n692), .C2(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n695), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT86), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G26), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n484), .A2(G128), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n482), .A2(G140), .ZN(new_n706));
  OR2_X1    g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  MUX2_X1   g286(.A(new_n704), .B(new_n711), .S(KEYINPUT28), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G2067), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n628), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G4), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(new_n715), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n719), .A2(KEYINPUT23), .A3(G20), .ZN(new_n720));
  AOI21_X1  g295(.A(KEYINPUT23), .B1(new_n719), .B2(G20), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n720), .B(new_n721), .C1(G299), .C2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1956), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n718), .B(new_n723), .C1(G2067), .C2(new_n712), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n530), .B2(new_n533), .ZN(new_n725));
  NOR2_X1   g300(.A1(G16), .A2(G22), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n725), .A2(G1971), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(G1971), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT33), .B(G1976), .Z(new_n730));
  AND3_X1   g305(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G16), .ZN(new_n732));
  OR2_X1    g307(.A1(G16), .A2(G23), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n719), .A2(G6), .ZN(new_n736));
  INV_X1    g311(.A(G305), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n719), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT32), .B(G1981), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n732), .A2(new_n733), .A3(new_n730), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n729), .A2(new_n735), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT91), .B1(new_n742), .B2(KEYINPUT34), .ZN(new_n743));
  INV_X1    g318(.A(new_n741), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(new_n734), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n745), .A2(new_n746), .A3(new_n729), .A4(new_n740), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n719), .A2(G24), .ZN(new_n748));
  INV_X1    g323(.A(G290), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n719), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT89), .B(G1986), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n750), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n703), .A2(G25), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n484), .A2(G119), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n482), .A2(G131), .ZN(new_n756));
  OR2_X1    g331(.A1(G95), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n703), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT35), .B(G1991), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT87), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT88), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n761), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n743), .A2(new_n747), .A3(new_n753), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n724), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n769), .A2(new_n770), .A3(new_n747), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n771), .A2(KEYINPUT36), .A3(new_n753), .A4(new_n765), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n703), .A2(G35), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n773), .B(new_n774), .C1(new_n486), .C2(G29), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT29), .B(G2090), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n768), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n780));
  AND3_X1   g355(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n482), .A2(G139), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n465), .A2(new_n467), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n784), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n475), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT94), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT92), .B1(G29), .B2(G33), .ZN(new_n789));
  OR3_X1    g364(.A1(KEYINPUT92), .A2(G29), .A3(G33), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT95), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n788), .A2(new_n793), .A3(new_n789), .A4(new_n790), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n792), .A2(G2072), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(G2072), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  OR2_X1    g371(.A1(G29), .A2(G32), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n482), .A2(G141), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT96), .Z(new_n799));
  AND3_X1   g374(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT26), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n800), .B(new_n802), .C1(G129), .C2(new_n484), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n797), .B1(new_n804), .B2(new_n703), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT27), .B(G1996), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n703), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n703), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n805), .A2(new_n806), .B1(new_n808), .B2(G2078), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT97), .B1(G5), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(KEYINPUT97), .A2(G5), .A3(G16), .ZN(new_n812));
  AOI211_X1 g387(.A(new_n811), .B(new_n812), .C1(G171), .C2(G16), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n809), .B1(G1961), .B2(new_n813), .C1(new_n805), .C2(new_n806), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n808), .A2(G2078), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n795), .A2(new_n796), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G34), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT24), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(KEYINPUT24), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n703), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G160), .B2(new_n703), .ZN(new_n821));
  INV_X1    g396(.A(G2084), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n813), .A2(G1961), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT98), .Z(new_n825));
  NOR2_X1   g400(.A1(G16), .A2(G21), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G168), .B2(G16), .ZN(new_n827));
  INV_X1    g402(.A(G1966), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n653), .A2(new_n703), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT31), .B(G11), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(G28), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(G28), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n834), .A3(new_n703), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n825), .A2(new_n836), .A3(KEYINPUT99), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n816), .B(new_n823), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n719), .A2(G19), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n557), .B2(new_n719), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(G1341), .Z(new_n847));
  NAND4_X1  g422(.A1(new_n779), .A2(new_n843), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n841), .B(KEYINPUT100), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n768), .A2(new_n772), .A3(new_n847), .A4(new_n778), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT102), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(G311));
  NAND3_X1  g427(.A1(new_n779), .A2(new_n843), .A3(new_n847), .ZN(G150));
  AOI22_X1  g428(.A1(new_n537), .A2(G55), .B1(new_n539), .B2(G93), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n513), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NOR2_X1   g433(.A1(new_n627), .A2(new_n635), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT39), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n856), .B(new_n557), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  OAI21_X1  g439(.A(new_n858), .B1(new_n864), .B2(G860), .ZN(G145));
  XNOR2_X1  g440(.A(new_n501), .B(new_n709), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n804), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(KEYINPUT104), .A3(new_n787), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n787), .A2(KEYINPUT104), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n787), .A2(KEYINPUT104), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n871), .B2(new_n867), .ZN(new_n872));
  AOI22_X1  g447(.A1(G130), .A2(new_n484), .B1(new_n482), .B2(G142), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n875), .B(new_n876), .C1(G118), .C2(new_n475), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n647), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n872), .A2(new_n879), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n653), .B(new_n477), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n486), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n760), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n880), .B2(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  AND3_X1   g464(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n590), .B1(new_n585), .B2(new_n589), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n890), .A2(new_n891), .A3(new_n627), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n625), .B1(new_n584), .B2(G92), .ZN(new_n893));
  INV_X1    g468(.A(G92), .ZN(new_n894));
  AOI211_X1 g469(.A(KEYINPUT10), .B(new_n894), .C1(new_n582), .C2(new_n583), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n581), .A2(new_n591), .B1(new_n896), .B2(new_n624), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT41), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n628), .A2(new_n581), .A3(new_n591), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n627), .B1(new_n890), .B2(new_n891), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n637), .B(new_n863), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n899), .A2(new_n900), .A3(new_n905), .A4(new_n901), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n904), .A2(new_n897), .A3(new_n892), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n903), .A2(new_n910), .A3(new_n904), .A4(new_n906), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G288), .B(G290), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n530), .A2(new_n533), .A3(G305), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n737), .B1(new_n531), .B2(new_n534), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G288), .B(new_n749), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n916), .A2(new_n919), .B1(new_n922), .B2(KEYINPUT42), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n912), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n908), .A2(new_n924), .A3(new_n909), .A4(new_n911), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(G868), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT109), .B1(new_n856), .B2(new_n616), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n926), .A2(KEYINPUT109), .A3(G868), .A4(new_n927), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(G295));
  AND3_X1   g507(.A1(new_n930), .A2(KEYINPUT110), .A3(new_n931), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT110), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(G331));
  XNOR2_X1  g510(.A(G171), .B(G286), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n863), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n863), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n903), .A2(new_n906), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n916), .A2(new_n919), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n937), .A2(new_n900), .A3(new_n899), .A4(new_n938), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n886), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n898), .A2(new_n902), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n939), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n939), .A3(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n942), .B(KEYINPUT112), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n886), .B(new_n943), .C1(new_n954), .C2(new_n941), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n946), .B1(new_n955), .B2(KEYINPUT43), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n944), .B2(new_n945), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  MUX2_X1   g534(.A(new_n956), .B(new_n959), .S(KEYINPUT44), .Z(G397));
  INV_X1    g535(.A(new_n804), .ZN(new_n961));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n709), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n804), .A2(G1996), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n759), .A2(new_n763), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n968), .A2(new_n969), .B1(new_n964), .B2(new_n710), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n498), .A2(G2105), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n499), .A2(new_n491), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n784), .A2(new_n492), .A3(new_n490), .ZN(new_n975));
  AOI21_X1  g550(.A(G2105), .B1(new_n975), .B2(new_n488), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n970), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n961), .B2(new_n965), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n982), .A2(KEYINPUT46), .A3(new_n962), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n982), .B2(new_n962), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  INV_X1    g564(.A(new_n763), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n968), .B1(new_n760), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n982), .B1(new_n991), .B2(new_n969), .ZN(new_n992));
  OR2_X1    g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n983), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT48), .Z(new_n995));
  AOI211_X1 g570(.A(new_n984), .B(new_n989), .C1(new_n992), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n495), .B2(new_n500), .ZN(new_n997));
  INV_X1    g572(.A(new_n981), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT119), .B(G8), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G305), .A2(G1981), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n539), .A2(G86), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n608), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1003), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1002), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n731), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1002), .B1(new_n1013), .B2(new_n1004), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n501), .A2(new_n971), .A3(new_n978), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n998), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n997), .A2(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n828), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n981), .B1(new_n997), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n822), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(G168), .A3(new_n1000), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1001), .B1(new_n731), .B2(G1976), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(new_n1027), .C1(G1976), .C2(new_n731), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1011), .B(new_n1028), .C1(new_n1027), .C2(new_n1026), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n980), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n981), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n977), .A2(KEYINPUT114), .A3(new_n979), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1031), .A2(KEYINPUT115), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1971), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G2090), .ZN(new_n1040));
  OR3_X1    g615(.A1(new_n1038), .A2(KEYINPUT117), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(G8), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(KEYINPUT118), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(KEYINPUT118), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1025), .B(new_n1029), .C1(new_n1043), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1014), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT56), .B(G2072), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1034), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n471), .A2(new_n476), .A3(G40), .A4(new_n1020), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n999), .A2(KEYINPUT121), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n998), .C1(new_n997), .C2(new_n1020), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n997), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1956), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT122), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1055), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n573), .A2(new_n580), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n585), .A2(new_n589), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(KEYINPUT123), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1069), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(KEYINPUT123), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(KEYINPUT57), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n999), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1039), .A2(new_n716), .B1(new_n964), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1068), .B2(new_n1079), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1080), .B1(new_n1083), .B2(new_n628), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1055), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1062), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1066), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT61), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n627), .A2(KEYINPUT126), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1082), .B2(KEYINPUT60), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n627), .A2(KEYINPUT126), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1082), .A2(new_n1095), .A3(KEYINPUT60), .A4(new_n1091), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT124), .B(G1996), .Z(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT58), .B(G1341), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1034), .A2(new_n1097), .B1(new_n1081), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n557), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1094), .A2(new_n1096), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1102), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1099), .A2(new_n557), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1079), .A4(new_n1085), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1090), .A2(new_n1103), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1084), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G2078), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1036), .A2(new_n1112), .A3(new_n1037), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n998), .B1(new_n977), .B2(new_n1019), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n997), .A2(new_n1060), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G1961), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1032), .A2(new_n980), .A3(KEYINPUT53), .A4(new_n1112), .ZN(new_n1121));
  XNOR2_X1  g696(.A(G171), .B(KEYINPUT54), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1115), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G8), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G286), .A2(new_n1000), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT51), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1015), .B(new_n998), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1118), .A2(new_n822), .B1(new_n1132), .B2(new_n828), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1000), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1133), .A2(new_n1126), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1132), .A2(new_n1114), .A3(G2078), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1119), .B(new_n1140), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1123), .B(new_n1139), .C1(new_n1141), .C2(new_n1122), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1052), .B1(new_n1111), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1025), .A2(KEYINPUT63), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1130), .B1(new_n1024), .B2(new_n1000), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1126), .B1(new_n1133), .B2(new_n1124), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(KEYINPUT51), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1146), .B(KEYINPUT62), .C1(new_n1149), .C2(new_n1137), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1137), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT127), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1139), .A2(KEYINPUT62), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1156));
  OAI21_X1  g731(.A(G171), .B1(new_n1156), .B2(new_n1140), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1145), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1029), .B1(new_n1144), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1062), .A2(G2090), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1000), .B1(new_n1038), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1048), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1051), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n969), .B(new_n991), .C1(G1986), .C2(G290), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n983), .B1(new_n1165), .B2(new_n993), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n996), .B1(new_n1164), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g742(.A1(G401), .A2(new_n461), .A3(G229), .ZN(new_n1169));
  INV_X1    g743(.A(G227), .ZN(new_n1170));
  NAND4_X1  g744(.A1(new_n956), .A2(new_n1169), .A3(new_n1170), .A4(new_n888), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


