//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G50), .B2(G226), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR3_X1   g0029(.A1(new_n221), .A2(new_n226), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n224), .A3(G1), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G58), .A2(G68), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n224), .B1(new_n222), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT7), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n255), .B1(new_n260), .B2(G20), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n254), .B1(new_n266), .B2(G68), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G159), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT16), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n267), .A2(new_n275), .A3(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n225), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n252), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n260), .B1(G226), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G223), .A2(G1698), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n282), .A2(new_n283), .B1(new_n257), .B2(new_n209), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT67), .ZN(new_n290));
  INV_X1    g0090(.A(new_n285), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G232), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT66), .B(G45), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(G274), .C1(new_n294), .C2(G41), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT72), .B1(new_n292), .B2(new_n295), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n286), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(new_n279), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G1), .B2(new_n224), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(new_n247), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n280), .A2(new_n300), .A3(new_n301), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT17), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n267), .A2(new_n275), .A3(new_n272), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n275), .B1(new_n267), .B2(new_n272), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n279), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n252), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(new_n304), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n298), .A2(G179), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n298), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT18), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n260), .B1(G232), .B2(new_n281), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G226), .A2(G1698), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n285), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT71), .ZN(new_n324));
  INV_X1    g0124(.A(new_n295), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n290), .A2(new_n291), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(G238), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(G179), .A3(new_n331), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT14), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n336), .A3(G169), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n224), .A2(G33), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n269), .A2(new_n202), .B1(new_n339), .B2(new_n217), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n224), .A2(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n279), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  INV_X1    g0143(.A(G68), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n342), .A2(new_n343), .B1(new_n344), .B2(new_n303), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n342), .A2(new_n343), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(new_n293), .A3(G13), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n347), .B(KEYINPUT12), .Z(new_n348));
  NOR3_X1   g0148(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n338), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n332), .B2(new_n299), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n329), .B2(new_n331), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  INV_X1    g0157(.A(new_n339), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n248), .A2(new_n268), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n224), .B2(new_n217), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n279), .B1(new_n217), .B2(new_n250), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n217), .B2(new_n303), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n325), .B1(new_n326), .B2(G244), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n264), .B1(G232), .B2(new_n281), .ZN(new_n365));
  INV_X1    g0165(.A(G238), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n281), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G107), .B2(new_n260), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n364), .B1(new_n291), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G200), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n363), .B(new_n370), .C1(new_n299), .C2(new_n369), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n318), .A2(new_n351), .A3(new_n356), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n250), .A2(G50), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n303), .B2(G50), .ZN(new_n374));
  XOR2_X1   g0174(.A(new_n374), .B(KEYINPUT68), .Z(new_n375));
  AOI22_X1  g0175(.A1(new_n248), .A2(new_n358), .B1(G20), .B2(new_n203), .ZN(new_n376));
  INV_X1    g0176(.A(G150), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n269), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n279), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT9), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n325), .B1(new_n326), .B2(G226), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n264), .B1(G222), .B2(new_n281), .ZN(new_n383));
  INV_X1    g0183(.A(G223), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n281), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(G77), .B2(new_n260), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n291), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G200), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n381), .B(new_n388), .C1(new_n299), .C2(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT70), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT10), .ZN(new_n391));
  OR3_X1    g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n387), .A2(G179), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n387), .A2(new_n314), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n380), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n369), .A2(G179), .ZN(new_n400));
  XOR2_X1   g0200(.A(new_n400), .B(KEYINPUT69), .Z(new_n401));
  NAND2_X1  g0201(.A1(new_n369), .A2(new_n314), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n362), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n372), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n293), .A2(G45), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT74), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n288), .A2(G1), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G41), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT75), .ZN(new_n415));
  INV_X1    g0215(.A(G274), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(KEYINPUT5), .B2(new_n287), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n408), .A2(new_n418), .A3(new_n413), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n415), .A2(new_n291), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(G250), .B(new_n281), .C1(new_n262), .C2(new_n263), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT86), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT86), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n260), .A2(new_n423), .A3(G250), .A4(new_n281), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G294), .ZN(new_n426));
  OAI211_X1 g0226(.A(G257), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT87), .ZN(new_n429));
  INV_X1    g0229(.A(new_n427), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n422), .B2(new_n424), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT87), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n426), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n291), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n420), .B1(new_n434), .B2(KEYINPUT88), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n431), .A2(new_n432), .A3(new_n426), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n431), .B2(new_n426), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT88), .B(new_n285), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n408), .A2(new_n439), .A3(new_n413), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G264), .A3(new_n291), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT89), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n420), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n285), .B1(new_n436), .B2(new_n437), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT88), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n441), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n434), .B2(KEYINPUT88), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT89), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n443), .A2(new_n451), .A3(new_n299), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n434), .A2(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n420), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n353), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n250), .A2(new_n279), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n293), .A2(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n251), .A2(G107), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(G20), .B1(new_n258), .B2(new_n259), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G87), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT22), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n224), .A2(G107), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT23), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(new_n470), .C1(G20), .C2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT24), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n461), .B(new_n465), .C1(new_n473), .C2(new_n279), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n456), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n314), .B1(new_n443), .B2(new_n451), .ZN(new_n476));
  INV_X1    g0276(.A(G179), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n454), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n279), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n460), .B2(new_n459), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n476), .A2(new_n478), .B1(new_n480), .B2(new_n465), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n250), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n224), .C1(G33), .C2(new_n211), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n279), .C1(new_n224), .C2(G116), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT20), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  OAI221_X1 g0290(.A(new_n484), .B1(new_n483), .B2(new_n459), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G264), .A2(G1698), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n260), .B(new_n492), .C1(new_n212), .C2(G1698), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n285), .C1(G303), .C2(new_n260), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n440), .A2(G270), .A3(new_n291), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n420), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n496), .A3(G169), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n498), .A2(KEYINPUT83), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n499), .ZN(new_n501));
  INV_X1    g0301(.A(new_n496), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(KEYINPUT82), .A3(G179), .A4(new_n491), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  INV_X1    g0304(.A(new_n491), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n420), .A2(G179), .A3(new_n494), .A4(new_n495), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n500), .A2(new_n501), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n505), .B1(new_n502), .B2(new_n353), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n509), .B(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n502), .A2(G190), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n440), .A2(G257), .A3(new_n291), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT76), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n440), .A2(KEYINPUT76), .A3(G257), .A4(new_n291), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n420), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT77), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n264), .A2(new_n218), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(KEYINPUT4), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(KEYINPUT4), .A3(new_n281), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n522), .A2(new_n523), .A3(new_n485), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT4), .B1(new_n264), .B2(new_n210), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n285), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n517), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n520), .A2(new_n477), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n251), .A2(G97), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n532));
  XOR2_X1   g0332(.A(G97), .B(G107), .Z(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(KEYINPUT6), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT73), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n268), .A2(G77), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(G20), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n266), .A2(G107), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n535), .C2(new_n536), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n531), .B1(new_n539), .B2(new_n279), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n211), .B2(new_n459), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n517), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT77), .B1(new_n517), .B2(new_n420), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n291), .B1(new_n524), .B2(new_n526), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n530), .B(new_n541), .C1(new_n545), .C2(G169), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n457), .A2(G97), .A3(new_n458), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n520), .A2(G190), .A3(new_n528), .A4(new_n529), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n545), .C2(new_n353), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n224), .A2(G33), .A3(G97), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT79), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n224), .B1(new_n319), .B2(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n209), .A2(new_n211), .A3(new_n460), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n224), .B(G68), .C1(new_n262), .C2(new_n263), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT80), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n551), .A2(new_n553), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT79), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n466), .A2(G68), .B1(new_n557), .B2(new_n558), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT80), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n569), .A3(new_n279), .ZN(new_n570));
  INV_X1    g0370(.A(new_n357), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n250), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT81), .B1(new_n459), .B2(new_n571), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT81), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n457), .A2(new_n574), .A3(new_n357), .A4(new_n458), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n570), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n218), .A2(G1698), .ZN(new_n578));
  OAI221_X1 g0378(.A(new_n578), .B1(G238), .B2(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n291), .B1(new_n579), .B2(new_n471), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n416), .B1(new_n210), .B2(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n409), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n407), .A2(KEYINPUT78), .A3(G250), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n285), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n314), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n477), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n577), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n579), .A2(new_n471), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n285), .ZN(new_n591));
  INV_X1    g0391(.A(new_n584), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n353), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n580), .A2(new_n299), .A3(new_n584), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n457), .A2(G87), .A3(new_n458), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n572), .A3(new_n570), .A4(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n546), .A2(new_n550), .A3(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n405), .A2(new_n482), .A3(new_n512), .A4(new_n599), .ZN(G372));
  INV_X1    g0400(.A(new_n398), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n355), .B(new_n307), .C1(new_n351), .C2(new_n403), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n602), .A2(new_n317), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n392), .A2(new_n395), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT90), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n589), .A2(new_n597), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n589), .B2(new_n597), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n609), .A2(new_n546), .A3(new_n550), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n435), .A2(new_n442), .A3(KEYINPUT89), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n450), .B1(new_n447), .B2(new_n449), .ZN(new_n612));
  OAI21_X1  g0412(.A(G169), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n478), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n474), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n610), .B(new_n475), .C1(new_n615), .C2(new_n508), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n607), .A2(new_n608), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n546), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT91), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n546), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .A3(new_n598), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT91), .B(new_n617), .C1(new_n618), .C2(new_n546), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n616), .A2(new_n625), .A3(new_n589), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n405), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n605), .A2(new_n627), .ZN(G369));
  NOR2_X1   g0428(.A1(new_n249), .A2(G20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n293), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n505), .A2(new_n636), .ZN(new_n637));
  MUX2_X1   g0437(.A(new_n512), .B(new_n508), .S(new_n637), .Z(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n475), .B(new_n481), .C1(new_n474), .C2(new_n636), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n481), .B2(new_n636), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n635), .B(KEYINPUT92), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n615), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n508), .A2(new_n636), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n482), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(G399));
  INV_X1    g0449(.A(new_n227), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G41), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n558), .A2(G116), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G1), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n223), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT26), .B1(new_n618), .B2(new_n546), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n589), .B(KEYINPUT95), .Z(new_n658));
  AOI21_X1  g0458(.A(new_n548), .B1(new_n545), .B2(new_n477), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n520), .A2(new_n528), .A3(new_n529), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n314), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(new_n617), .A3(new_n661), .A4(new_n598), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT96), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT96), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n657), .A2(new_n665), .A3(new_n658), .A4(new_n662), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n616), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n636), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT29), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n626), .A2(new_n645), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(KEYINPUT29), .B2(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n546), .A2(new_n550), .A3(new_n598), .A4(new_n645), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n475), .A2(new_n672), .A3(new_n481), .A4(new_n512), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n520), .A2(new_n528), .A3(new_n529), .A4(new_n585), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n506), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n506), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n675), .A2(new_n676), .A3(new_n453), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n453), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT30), .B1(new_n682), .B2(new_n674), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n502), .A2(G179), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n454), .A2(new_n660), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n586), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n681), .A2(new_n683), .B1(new_n686), .B2(new_n586), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n636), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n673), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT94), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(KEYINPUT94), .A3(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n671), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n656), .B1(new_n699), .B2(G1), .ZN(G364));
  XNOR2_X1  g0500(.A(new_n629), .B(KEYINPUT97), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n293), .B1(new_n701), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n651), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n650), .A2(new_n260), .ZN(new_n706));
  OAI221_X1 g0506(.A(new_n706), .B1(new_n223), .B2(new_n294), .C1(new_n242), .C2(new_n288), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n260), .A2(G355), .A3(new_n227), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n707), .B(new_n708), .C1(G116), .C2(new_n227), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n225), .B1(G20), .B2(new_n314), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n705), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n712), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n224), .A2(new_n299), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n477), .A2(G200), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n224), .A2(G190), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(G322), .A2(new_n719), .B1(new_n723), .B2(G329), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n353), .A2(G179), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n717), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G303), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n720), .A2(new_n725), .ZN(new_n732));
  INV_X1    g0532(.A(G283), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G190), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(KEYINPUT99), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(KEYINPUT99), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT33), .B(G317), .Z(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n224), .B1(new_n721), .B2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n260), .B1(new_n743), .B2(G294), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n735), .A2(new_n299), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G326), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n720), .A2(new_n718), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n744), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n731), .A2(new_n734), .A3(new_n741), .A4(new_n749), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n722), .A2(KEYINPUT32), .A3(new_n270), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n745), .A2(G50), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT32), .B1(new_n722), .B2(new_n270), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n743), .A2(G97), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n729), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G87), .ZN(new_n757));
  INV_X1    g0557(.A(new_n732), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n264), .B1(new_n758), .B2(G107), .ZN(new_n759));
  INV_X1    g0559(.A(G58), .ZN(new_n760));
  INV_X1    g0560(.A(new_n719), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n757), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n739), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n755), .B(new_n762), .C1(G68), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n748), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G77), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n750), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT100), .Z(new_n768));
  INV_X1    g0568(.A(new_n713), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n715), .B1(new_n638), .B2(new_n716), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n639), .A2(new_n705), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n638), .A2(G330), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(G396));
  NAND2_X1  g0573(.A1(new_n745), .A2(G303), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n754), .A2(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n260), .B(new_n775), .C1(G87), .C2(new_n758), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n761), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n739), .A2(new_n733), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G116), .A2(new_n765), .B1(new_n723), .B2(G311), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n729), .B2(new_n460), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n777), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n719), .A2(G143), .B1(G137), .B2(new_n745), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n784), .B1(new_n270), .B2(new_n748), .C1(new_n739), .C2(new_n377), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n758), .A2(G68), .ZN(new_n788));
  INV_X1    g0588(.A(G132), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n760), .B2(new_n742), .C1(new_n789), .C2(new_n722), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n264), .B1(new_n756), .B2(G50), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n783), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n713), .A2(new_n710), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n793), .A2(new_n769), .B1(G77), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n404), .A2(new_n636), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n371), .B1(new_n363), .B2(new_n636), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n403), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n705), .B(new_n796), .C1(new_n800), .C2(new_n710), .ZN(new_n801));
  INV_X1    g0601(.A(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n698), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n800), .B1(new_n696), .B2(new_n697), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(new_n670), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n801), .B1(new_n806), .B2(new_n705), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G384));
  INV_X1    g0608(.A(KEYINPUT38), .ZN(new_n809));
  INV_X1    g0609(.A(new_n633), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n312), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n305), .B(KEYINPUT17), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT18), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n316), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT102), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n305), .A2(new_n316), .A3(new_n811), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n818), .A2(new_n305), .A3(new_n316), .A4(new_n811), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n809), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n811), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n307), .B2(new_n317), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n826), .A2(KEYINPUT38), .A3(new_n821), .A4(new_n822), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(KEYINPUT39), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n351), .A2(new_n635), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n305), .A2(new_n316), .A3(KEYINPUT103), .A4(new_n811), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n816), .A3(new_n832), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n826), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n809), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(new_n827), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n828), .B(new_n829), .C1(new_n838), .C2(KEYINPUT39), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n317), .A2(new_n633), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n350), .A2(new_n635), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n351), .A2(new_n356), .A3(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n350), .B(new_n635), .C1(new_n338), .C2(new_n355), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n626), .A2(new_n645), .A3(new_n799), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n797), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n824), .A2(new_n827), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n839), .A2(new_n840), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n671), .A2(new_n405), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n605), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n849), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n842), .A2(new_n843), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n635), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n673), .A2(new_n854), .A3(new_n692), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n847), .A2(new_n802), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n837), .B2(new_n827), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n802), .A2(new_n855), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n844), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n405), .A2(new_n855), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G330), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n852), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n293), .B2(new_n701), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n483), .B1(new_n534), .B2(KEYINPUT35), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n225), .A2(new_n224), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n869), .B(new_n870), .C1(KEYINPUT35), .C2(new_n534), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT36), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n253), .A2(G77), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n223), .A2(new_n873), .B1(G50), .B2(new_n344), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(G1), .A3(new_n249), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n868), .A2(new_n872), .A3(new_n875), .ZN(G367));
  NAND2_X1  g0676(.A1(new_n622), .A2(new_n644), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n546), .B(new_n550), .C1(new_n548), .C2(new_n645), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n482), .A2(new_n647), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n546), .B1(new_n481), .B2(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n645), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(new_n887), .A3(new_n883), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT104), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n570), .A2(new_n572), .A3(new_n596), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n635), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n609), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n589), .B2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n890), .B1(new_n889), .B2(new_n895), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n896), .A2(new_n897), .B1(KEYINPUT43), .B2(new_n894), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n889), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT104), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n643), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n879), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n699), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n648), .A2(new_n646), .A3(new_n879), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT45), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n648), .A2(KEYINPUT45), .A3(new_n646), .A4(new_n879), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n648), .A2(new_n646), .ZN(new_n916));
  INV_X1    g0716(.A(new_n879), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT44), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT44), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(new_n643), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n648), .B1(new_n642), .B2(new_n647), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n639), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n910), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n651), .B(KEYINPUT41), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n702), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n898), .A2(new_n903), .A3(KEYINPUT106), .A4(new_n905), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n909), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n202), .A2(new_n748), .B1(new_n732), .B2(new_n217), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n756), .B2(G58), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n742), .A2(new_n344), .ZN(new_n935));
  INV_X1    g0735(.A(G137), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n260), .B1(new_n722), .B2(new_n936), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n935), .B(new_n937), .C1(G143), .C2(new_n745), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n939), .B1(new_n377), .B2(new_n761), .C1(new_n270), .C2(new_n739), .ZN(new_n940));
  INV_X1    g0740(.A(new_n745), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n264), .B1(new_n742), .B2(new_n460), .C1(new_n941), .C2(new_n747), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n723), .A2(G317), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(new_n211), .B2(new_n732), .C1(new_n761), .C2(new_n730), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(G283), .C2(new_n765), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n729), .A2(new_n483), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n946), .A2(KEYINPUT46), .B1(G294), .B2(new_n763), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n945), .B(new_n947), .C1(KEYINPUT46), .C2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n940), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n705), .B1(new_n950), .B2(new_n713), .ZN(new_n951));
  INV_X1    g0751(.A(new_n706), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n714), .B1(new_n227), .B2(new_n571), .C1(new_n237), .C2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n894), .C2(new_n716), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n932), .A2(new_n954), .ZN(G387));
  NAND2_X1  g0755(.A1(new_n910), .A2(new_n925), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n926), .A2(new_n699), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n957), .A3(new_n651), .ZN(new_n958));
  INV_X1    g0758(.A(new_n294), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n706), .B1(new_n234), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n653), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(new_n227), .A3(new_n260), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n344), .A2(new_n217), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n248), .A2(new_n202), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n961), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n966), .B(new_n288), .C1(KEYINPUT50), .C2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n963), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n650), .A2(new_n460), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n713), .B(new_n712), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n739), .A2(new_n247), .B1(new_n344), .B2(new_n748), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT107), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n260), .B1(new_n722), .B2(new_n377), .C1(new_n211), .C2(new_n732), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n571), .A2(new_n742), .B1(new_n270), .B2(new_n941), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n756), .C2(G77), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(new_n975), .C1(new_n202), .C2(new_n761), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT108), .Z(new_n977));
  AOI22_X1  g0777(.A1(new_n719), .A2(G317), .B1(G322), .B2(new_n745), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n730), .B2(new_n748), .C1(new_n739), .C2(new_n747), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT109), .Z(new_n980));
  AOI22_X1  g0780(.A1(new_n980), .A2(KEYINPUT48), .B1(G283), .B2(new_n743), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(KEYINPUT48), .B2(new_n980), .C1(new_n778), .C2(new_n729), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n260), .B1(new_n723), .B2(G326), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n732), .A2(new_n483), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n705), .B(new_n970), .C1(new_n989), .C2(new_n713), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(KEYINPUT111), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n642), .C2(new_n716), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n926), .A2(new_n703), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n958), .A2(new_n993), .A3(new_n994), .ZN(G393));
  INV_X1    g0795(.A(new_n957), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n923), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n922), .A2(new_n904), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT112), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n922), .A2(new_n904), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n922), .A2(new_n999), .A3(new_n904), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n997), .B(new_n651), .C1(new_n1003), .C2(new_n996), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n917), .A2(new_n712), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n714), .B1(new_n211), .B2(new_n227), .C1(new_n245), .C2(new_n952), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n264), .B1(new_n732), .B2(new_n460), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G322), .B2(new_n723), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n483), .B2(new_n742), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G283), .B2(new_n756), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n778), .B2(new_n748), .C1(new_n730), .C2(new_n739), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n719), .A2(G311), .B1(G317), .B2(new_n745), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT52), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n756), .A2(G68), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n763), .A2(G50), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n723), .A2(G143), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n260), .B1(new_n732), .B2(new_n209), .C1(new_n247), .C2(new_n748), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G77), .B2(new_n743), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n719), .A2(G159), .B1(G150), .B2(new_n745), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1011), .A2(new_n1013), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n705), .B1(new_n1023), .B2(new_n713), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1005), .A2(new_n1006), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1003), .B2(new_n703), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1004), .A2(new_n1026), .ZN(G390));
  NAND2_X1  g0827(.A1(new_n845), .A2(new_n797), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n853), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n829), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n828), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT115), .B1(new_n846), .B2(new_n829), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n667), .A2(new_n636), .A3(new_n799), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n797), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT114), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1039), .A3(new_n797), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n853), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n838), .A2(new_n829), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n693), .A2(KEYINPUT94), .A3(G330), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT94), .B1(new_n693), .B2(G330), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n802), .B(new_n853), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n1035), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(G330), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n860), .A2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1035), .A2(new_n1043), .B1(new_n853), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n703), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1033), .A2(new_n710), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n260), .B1(new_n745), .B2(G283), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n788), .B(new_n1054), .C1(new_n217), .C2(new_n742), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n757), .B1(new_n211), .B2(new_n748), .C1(new_n483), .C2(new_n761), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G107), .C2(new_n763), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n723), .A2(G294), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n260), .B1(new_n761), .B2(new_n789), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G50), .B2(new_n758), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n723), .A2(G125), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT54), .B(G143), .Z(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT117), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n765), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n743), .A2(G159), .B1(G128), .B2(new_n745), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G137), .B2(new_n763), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n729), .A2(new_n377), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT53), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1057), .A2(new_n1058), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n704), .B1(new_n248), .B2(new_n795), .C1(new_n1070), .C2(new_n769), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT118), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1053), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1052), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n844), .B1(new_n860), .B2(new_n1049), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1040), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1039), .B1(new_n1036), .B2(new_n797), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1046), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1050), .A2(new_n853), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n804), .B2(new_n853), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1028), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1084), .A2(KEYINPUT116), .A3(new_n1046), .A4(new_n1075), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1080), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n864), .A2(G330), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n850), .A2(new_n605), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n1081), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1035), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n652), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1074), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G378));
  NAND2_X1  g0900(.A1(new_n399), .A2(KEYINPUT119), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT119), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n392), .A2(new_n1102), .A3(new_n395), .A4(new_n398), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n380), .A2(new_n810), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1101), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n710), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n794), .A2(new_n202), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n745), .A2(G125), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1112), .B1(new_n377), .B2(new_n742), .C1(new_n761), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n756), .B2(new_n1063), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n789), .B2(new_n739), .C1(new_n936), .C2(new_n748), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT59), .Z(new_n1117));
  AOI21_X1  g0917(.A(G41), .B1(new_n723), .B2(G124), .ZN(new_n1118));
  AOI21_X1  g0918(.A(G33), .B1(new_n758), .B2(G159), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n202), .B1(new_n262), .B2(G41), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n357), .A2(new_n765), .B1(new_n719), .B2(G107), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n729), .B2(new_n217), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n264), .B1(new_n732), .B2(new_n760), .C1(new_n941), .C2(new_n483), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(G41), .A4(new_n935), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n211), .B2(new_n739), .C1(new_n733), .C2(new_n722), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT58), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1120), .A2(new_n1121), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n705), .B1(new_n1128), .B2(new_n713), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1110), .A2(new_n1111), .A3(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n857), .A2(new_n856), .B1(new_n859), .B2(new_n861), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1109), .B1(new_n1131), .B2(G330), .ZN(new_n1132));
  AND4_X1   g0932(.A1(G330), .A2(new_n858), .A3(new_n862), .A4(new_n1109), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n849), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1109), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n863), .B2(new_n1049), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n839), .A2(new_n840), .A3(new_n848), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(G330), .A3(new_n1109), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1139), .A3(KEYINPUT120), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT120), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n849), .B(new_n1141), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1130), .B1(new_n1143), .B2(new_n702), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1089), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT57), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1088), .B1(new_n1094), .B2(new_n1086), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT57), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n651), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1145), .B1(new_n1148), .B2(new_n1152), .ZN(G375));
  OAI22_X1  g0953(.A1(new_n729), .A2(new_n211), .B1(new_n730), .B2(new_n722), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT121), .Z(new_n1155));
  OAI22_X1  g0955(.A1(new_n571), .A2(new_n742), .B1(new_n778), .B2(new_n941), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n264), .B1(new_n217), .B2(new_n732), .C1(new_n761), .C2(new_n733), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n763), .C2(G116), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1155), .B(new_n1158), .C1(new_n460), .C2(new_n748), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT122), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n761), .A2(new_n936), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n748), .A2(new_n377), .B1(new_n722), .B2(new_n1113), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n756), .B2(G159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n763), .A2(new_n1063), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n941), .A2(new_n789), .B1(new_n732), .B2(new_n760), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n264), .B(new_n1165), .C1(G50), .C2(new_n743), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1160), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n705), .B1(new_n1168), .B2(new_n713), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n853), .B2(new_n711), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n344), .B2(new_n794), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1086), .B2(new_n703), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1080), .A2(new_n1083), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n928), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1090), .B2(new_n1174), .ZN(G381));
  INV_X1    g0975(.A(new_n1151), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n652), .B1(new_n1146), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1144), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1099), .ZN(new_n1181));
  OR4_X1    g0981(.A1(G384), .A2(new_n1181), .A3(G387), .A4(G390), .ZN(new_n1182));
  OR2_X1    g0982(.A1(G393), .A2(G396), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(G381), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1182), .A2(new_n1184), .ZN(G407));
  OAI221_X1 g0985(.A(G213), .B1(G343), .B2(new_n1181), .C1(new_n1182), .C2(new_n1184), .ZN(G409));
  NAND3_X1  g0986(.A1(new_n932), .A2(new_n954), .A3(G390), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(G393), .B(G396), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(G390), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(G387), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(KEYINPUT126), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT126), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n932), .A2(G390), .A3(new_n1193), .A4(new_n954), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT125), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1188), .B(new_n1196), .ZN(new_n1197));
  AOI221_X4 g0997(.A(KEYINPUT127), .B1(new_n1189), .B2(new_n1191), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT127), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT123), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n634), .A2(G213), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1146), .A2(new_n1147), .A3(new_n928), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1150), .A2(new_n703), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1099), .A2(new_n1206), .A3(new_n1130), .A4(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1205), .B(new_n1208), .C1(new_n1180), .C2(new_n1099), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1173), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1097), .B1(new_n1210), .B2(KEYINPUT60), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT60), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n651), .B1(new_n1173), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1172), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n807), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G384), .B(new_n1172), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1204), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1208), .A2(new_n1205), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G375), .A2(G378), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1217), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(KEYINPUT123), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT62), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT62), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT124), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n634), .A2(G213), .A3(G2897), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1215), .A2(KEYINPUT124), .A3(new_n1216), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1227), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT124), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1217), .B2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1209), .A2(new_n1226), .A3(new_n1228), .A4(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1224), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1203), .B1(new_n1223), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1225), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1231), .A2(new_n1228), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT61), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT63), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1218), .A2(new_n1222), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1219), .A2(KEYINPUT63), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1235), .A2(new_n1243), .ZN(G405));
  NAND2_X1  g1044(.A1(new_n1220), .A2(new_n1181), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(new_n1221), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(new_n1241), .ZN(G402));
endmodule


