//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT31), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G113), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n191), .B(new_n193), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n193), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT2), .B(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  OAI21_X1  g023(.A(G128), .B1(new_n203), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n210), .B(new_n211), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n217), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n204), .B2(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n211), .B1(new_n221), .B2(new_n210), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT65), .B(new_n224), .C1(new_n225), .C2(G137), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G131), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(G137), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n229), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT65), .B1(new_n238), .B2(new_n224), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n236), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n237), .ZN(new_n247));
  AND2_X1   g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n221), .A2(new_n250), .B1(new_n205), .B2(new_n248), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n223), .A2(new_n242), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n201), .B1(new_n252), .B2(KEYINPUT30), .ZN(new_n253));
  AOI211_X1 g067(.A(G131), .B(new_n235), .C1(new_n228), .C2(new_n229), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n231), .B1(new_n230), .B2(new_n236), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n216), .A2(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n212), .A2(new_n214), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(new_n216), .ZN(new_n259));
  INV_X1    g073(.A(new_n207), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n217), .B1(new_n258), .B2(new_n216), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n206), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT66), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n264), .B2(new_n218), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n256), .B(KEYINPUT30), .C1(new_n265), .C2(new_n241), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n223), .A2(new_n242), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(KEYINPUT67), .A3(KEYINPUT30), .A4(new_n256), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n253), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n201), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n256), .B(new_n272), .C1(new_n265), .C2(new_n241), .ZN(new_n273));
  NOR2_X1   g087(.A1(G237), .A2(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G210), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT27), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G101), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n189), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n268), .A2(new_n270), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n256), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n272), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n279), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(KEYINPUT31), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n273), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n272), .B1(new_n269), .B2(new_n256), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT28), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n273), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n278), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n188), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n299));
  INV_X1    g113(.A(new_n278), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(new_n291), .A3(new_n299), .A4(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n291), .A2(new_n293), .A3(new_n278), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n301), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n278), .B1(new_n285), .B2(new_n273), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n297), .B(new_n303), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n296), .A2(KEYINPUT32), .B1(G472), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT31), .B1(new_n285), .B2(new_n286), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n189), .B(new_n279), .C1(new_n281), .C2(new_n284), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n295), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n187), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT68), .B(KEYINPUT32), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT69), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n316), .B(new_n313), .C1(new_n311), .C2(new_n187), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n308), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(G234), .B2(new_n297), .ZN(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT75), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G125), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n328), .A3(KEYINPUT73), .A4(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n216), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n333), .A2(new_n337), .A3(new_n340), .A4(G146), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n206), .A2(G119), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n190), .A2(G128), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n345), .B1(new_n351), .B2(new_n346), .ZN(new_n352));
  OAI21_X1  g166(.A(G110), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n345), .A2(new_n348), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT24), .B(G110), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n344), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n360));
  OAI211_X1 g174(.A(G119), .B(new_n206), .C1(new_n360), .C2(new_n350), .ZN(new_n361));
  INV_X1    g175(.A(G110), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n348), .A4(new_n347), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n355), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n338), .A2(new_n216), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n343), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n326), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n357), .B1(new_n342), .B2(new_n343), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n365), .A2(new_n343), .A3(new_n366), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT74), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n325), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n325), .B1(new_n359), .B2(new_n367), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n375), .B2(new_n297), .ZN(new_n376));
  INV_X1    g190(.A(new_n325), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n359), .A2(new_n326), .A3(new_n367), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT74), .B1(new_n369), .B2(new_n370), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT25), .B(new_n297), .C1(new_n380), .C2(new_n373), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n320), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n320), .A2(G902), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT76), .Z(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  INV_X1    g206(.A(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n391), .A2(new_n394), .A3(new_n398), .A4(new_n395), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n401), .A3(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n201), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n404));
  INV_X1    g218(.A(new_n395), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n390), .A2(G107), .ZN(new_n406));
  OAI21_X1  g220(.A(G101), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n399), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT5), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n410), .B(G113), .C1(KEYINPUT5), .C2(new_n191), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n197), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n400), .A2(new_n413), .A3(new_n201), .A4(new_n402), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G122), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n404), .A2(new_n412), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n416), .A2(KEYINPUT6), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n412), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n201), .A2(new_n402), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n413), .B1(new_n420), .B2(new_n400), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n412), .A4(new_n414), .ZN(new_n423));
  INV_X1    g237(.A(new_n415), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n265), .A2(new_n334), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n251), .A2(new_n334), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G224), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n422), .A2(new_n423), .A3(new_n433), .A4(new_n424), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n426), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n431), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n427), .A2(KEYINPUT7), .A3(new_n428), .A4(new_n436), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n415), .B(KEYINPUT81), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT8), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n411), .A2(new_n197), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n408), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n412), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n438), .A2(new_n416), .A3(new_n439), .A4(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(new_n297), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n435), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT82), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n450), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n435), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n251), .A2(new_n400), .A3(new_n402), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n209), .B1(new_n258), .B2(new_n216), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n259), .B1(new_n458), .B2(new_n206), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n408), .B1(new_n459), .B2(new_n208), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(KEYINPUT10), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n409), .A2(KEYINPUT10), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n265), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n247), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n409), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n205), .B1(G128), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n409), .B1(new_n467), .B2(new_n261), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT77), .B1(new_n254), .B2(new_n255), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT77), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n246), .A2(new_n472), .A3(new_n237), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n465), .A2(new_n470), .A3(new_n474), .A4(new_n457), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n464), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n321), .A2(G227), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n479), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n254), .A2(new_n255), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n208), .B(new_n408), .C1(new_n219), .C2(new_n222), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n468), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n487));
  AOI211_X1 g301(.A(new_n487), .B(new_n482), .C1(new_n483), .C2(new_n468), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n475), .B(new_n481), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n297), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n475), .B1(new_n486), .B2(new_n488), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n479), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n461), .A2(new_n463), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n479), .B1(new_n495), .B2(new_n474), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n464), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(G469), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n491), .A2(new_n297), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT9), .B(G234), .ZN(new_n502));
  OAI21_X1  g316(.A(G221), .B1(new_n502), .B2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n390), .ZN(new_n506));
  INV_X1    g320(.A(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n321), .A3(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT84), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n274), .A2(new_n510), .A3(G214), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n204), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n509), .A2(KEYINPUT85), .A3(new_n204), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n507), .A2(new_n321), .A3(G143), .A4(G214), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n231), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT18), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n519), .B1(new_n514), .B2(new_n515), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n338), .A2(new_n216), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n523), .A2(new_n524), .B1(new_n366), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  AOI211_X1 g341(.A(G131), .B(new_n519), .C1(new_n514), .C2(new_n515), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n528), .A2(new_n521), .A3(KEYINPUT17), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n510), .B1(new_n274), .B2(G214), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(new_n258), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT85), .B1(new_n531), .B2(new_n511), .ZN(new_n532));
  INV_X1    g346(.A(new_n515), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n520), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT17), .A3(G131), .ZN(new_n535));
  INV_X1    g349(.A(new_n344), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n506), .B(new_n527), .C1(new_n529), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n506), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n523), .A2(new_n524), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n525), .A2(new_n366), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n523), .A2(new_n543), .A3(new_n231), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n338), .B1(KEYINPUT87), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n547), .B(new_n216), .C1(new_n338), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n343), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n534), .A2(G131), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n523), .A2(new_n231), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n539), .B1(new_n545), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n538), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NOR2_X1   g370(.A1(G475), .A2(G902), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT88), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n538), .B2(new_n554), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g379(.A(G122), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G116), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n192), .A2(G122), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n569), .B1(new_n567), .B2(new_n568), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n393), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n206), .A2(G143), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n258), .B2(new_n206), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G134), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n225), .B(new_n575), .C1(new_n258), .C2(new_n206), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n567), .A2(new_n568), .ZN(new_n581));
  OAI211_X1 g395(.A(G107), .B(new_n580), .C1(new_n581), .C2(KEYINPUT14), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n583), .B(new_n393), .C1(new_n571), .C2(new_n572), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n574), .A2(new_n579), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n204), .A2(new_n586), .A3(G128), .ZN(new_n587));
  OAI211_X1 g401(.A(G134), .B(new_n587), .C1(new_n576), .C2(new_n586), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n571), .A2(new_n393), .A3(new_n572), .ZN(new_n589));
  INV_X1    g403(.A(new_n572), .ZN(new_n590));
  AOI21_X1  g404(.A(G107), .B1(new_n590), .B2(new_n570), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n588), .B(new_n578), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n502), .A2(new_n319), .A3(G953), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n585), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n593), .B1(new_n585), .B2(new_n592), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n297), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n585), .A2(new_n592), .ZN(new_n600));
  INV_X1    g414(.A(new_n593), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n594), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT92), .A3(new_n297), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n565), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n604), .A2(new_n565), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n538), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT17), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n551), .A2(new_n609), .A3(new_n552), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n344), .B1(new_n521), .B2(KEYINPUT17), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n506), .B1(new_n612), .B2(new_n527), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n297), .B1(new_n608), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G475), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n321), .A2(G952), .ZN(new_n616));
  NAND2_X1  g430(.A1(G234), .A2(G237), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(G902), .A3(G953), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT21), .B(G898), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n563), .A2(new_n607), .A3(new_n615), .A4(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n456), .A2(new_n504), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n318), .A2(new_n389), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  AOI21_X1  g442(.A(new_n294), .B1(new_n280), .B2(new_n287), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT93), .B(G472), .C1(new_n629), .C2(G902), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT93), .ZN(new_n631));
  INV_X1    g445(.A(G472), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n311), .B(new_n297), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n455), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n451), .B2(new_n453), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n504), .A2(new_n388), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n603), .A2(KEYINPUT33), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n602), .A2(new_n640), .A3(new_n594), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(G478), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n603), .A2(new_n564), .A3(new_n297), .ZN(new_n643));
  NAND2_X1  g457(.A1(G478), .A2(G902), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n623), .B(new_n645), .C1(new_n563), .C2(new_n615), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n635), .A2(new_n637), .A3(new_n638), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT94), .Z(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT34), .B(G104), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n562), .A2(new_n561), .ZN(new_n652));
  INV_X1    g466(.A(new_n561), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n653), .B(new_n558), .C1(new_n538), .C2(new_n554), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n651), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n550), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n528), .B2(new_n521), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n506), .B1(new_n527), .B2(new_n657), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n610), .A2(new_n611), .B1(new_n522), .B2(new_n526), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n506), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n653), .B1(new_n660), .B2(new_n558), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n562), .A2(new_n561), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(KEYINPUT95), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n605), .ZN(new_n665));
  INV_X1    g479(.A(new_n606), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n665), .A2(new_n666), .B1(new_n614), .B2(G475), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n623), .B(KEYINPUT96), .Z(new_n669));
  NAND3_X1  g483(.A1(new_n454), .A2(new_n455), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n635), .A3(new_n638), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n378), .A2(new_n379), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n675), .A2(KEYINPUT36), .A3(new_n325), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n675), .B1(KEYINPUT36), .B2(new_n325), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n385), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n383), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n630), .A2(new_n633), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT97), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT97), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n630), .A2(new_n633), .A3(new_n683), .A4(new_n680), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n626), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  INV_X1    g501(.A(KEYINPUT98), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT25), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n373), .B1(new_n675), .B2(new_n325), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(G902), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n381), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n678), .B1(new_n692), .B2(new_n320), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n504), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n615), .B1(new_n605), .B2(new_n606), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n655), .B2(new_n663), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n620), .A2(G900), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n618), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n694), .A2(new_n696), .A3(new_n637), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n305), .A2(new_n306), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n303), .A2(new_n297), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n311), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n316), .B1(new_n296), .B2(new_n313), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n312), .A2(KEYINPUT69), .A3(new_n314), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n688), .B1(new_n699), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n503), .ZN(new_n709));
  AOI21_X1  g523(.A(G902), .B1(new_n480), .B2(new_n489), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n499), .B1(new_n710), .B2(new_n491), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n711), .B2(new_n498), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n637), .A2(new_n712), .A3(new_n680), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n652), .A2(new_n654), .A3(new_n651), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT95), .B1(new_n661), .B2(new_n662), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n667), .B(new_n698), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n318), .A3(KEYINPUT98), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n708), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G128), .ZN(G30));
  AND2_X1   g534(.A1(new_n451), .A2(new_n453), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT38), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n698), .B(KEYINPUT39), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n712), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n722), .B1(KEYINPUT40), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n285), .A2(new_n273), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n278), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n289), .A2(new_n290), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n728), .B2(new_n300), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n632), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n315), .B2(new_n317), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n724), .A2(KEYINPUT40), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n563), .A2(new_n615), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n636), .B1(new_n665), .B2(new_n666), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n693), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n725), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n258), .ZN(G45));
  INV_X1    g553(.A(new_n645), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n734), .A2(new_n740), .A3(new_n698), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n713), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n318), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G146), .ZN(G48));
  INV_X1    g558(.A(new_n487), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n484), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n484), .B2(new_n485), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n747), .A2(new_n496), .B1(new_n476), .B2(new_n479), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n748), .B2(G902), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n503), .A3(new_n492), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT99), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n749), .A2(new_n492), .A3(KEYINPUT99), .A4(new_n503), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n752), .A2(new_n637), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n318), .A2(new_n389), .A3(new_n646), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT100), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n755), .B(new_n757), .ZN(G15));
  AND2_X1   g572(.A1(new_n752), .A2(new_n753), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n318), .A2(new_n671), .A3(new_n389), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  NOR2_X1   g575(.A1(new_n625), .A2(new_n693), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n318), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  AND4_X1   g578(.A1(new_n454), .A2(new_n734), .A3(new_n735), .A4(new_n669), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n632), .B1(new_n311), .B2(new_n297), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n298), .A2(new_n291), .A3(new_n299), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n300), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n188), .B1(new_n288), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n766), .A2(new_n388), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  INV_X1    g586(.A(new_n741), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n766), .A2(new_n693), .A3(new_n769), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n754), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT101), .B(G125), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G27));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT32), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n629), .A2(new_n779), .A3(new_n188), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT32), .B1(new_n311), .B2(new_n187), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n629), .B2(new_n188), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT103), .A3(new_n703), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n702), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT102), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n498), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n494), .A2(KEYINPUT102), .A3(G469), .A4(new_n497), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n711), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n709), .A2(new_n636), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n721), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n741), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n389), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT42), .ZN(new_n794));
  INV_X1    g608(.A(new_n791), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n318), .A2(new_n389), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G131), .ZN(G33));
  INV_X1    g613(.A(new_n716), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n318), .A2(new_n800), .A3(new_n389), .A4(new_n795), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n563), .A2(new_n740), .A3(new_n615), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT43), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n634), .A2(new_n680), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n454), .A2(new_n636), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n805), .A2(new_n806), .A3(new_n803), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n494), .A2(new_n497), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(KEYINPUT45), .ZN(new_n813));
  OAI21_X1  g627(.A(G469), .B1(new_n812), .B2(KEYINPUT45), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT46), .B(new_n500), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(KEYINPUT104), .A3(new_n492), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT46), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n814), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(new_n499), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT104), .B1(new_n815), .B2(new_n492), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n503), .B(new_n723), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT105), .ZN(new_n823));
  INV_X1    g637(.A(new_n821), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n819), .A3(new_n816), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT105), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n503), .A4(new_n723), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT106), .B(G137), .Z(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(G39));
  INV_X1    g644(.A(KEYINPUT47), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n831), .A3(new_n503), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n503), .B1(new_n820), .B2(new_n821), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT47), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT108), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n773), .A2(new_n388), .A3(new_n808), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n318), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT107), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n834), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT108), .B1(new_n843), .B2(new_n840), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G140), .ZN(G42));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n698), .A2(new_n503), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n789), .A2(new_n693), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n454), .A2(new_n734), .A3(new_n735), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n318), .A2(new_n742), .B1(new_n732), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n717), .A2(new_n318), .A3(KEYINPUT98), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT98), .B1(new_n717), .B2(new_n318), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n852), .B(new_n775), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT52), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n760), .A2(new_n755), .A3(new_n763), .A4(new_n771), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n734), .A2(new_n740), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n670), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n635), .A2(new_n638), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n627), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n627), .A2(KEYINPUT110), .A3(new_n861), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n857), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n607), .A2(new_n615), .A3(new_n698), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n664), .A3(new_n712), .A4(new_n680), .ZN(new_n868));
  INV_X1    g682(.A(new_n808), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n870), .A2(new_n318), .B1(new_n792), .B2(new_n774), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n794), .A2(new_n797), .A3(new_n801), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n734), .A2(new_n607), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n635), .A2(new_n638), .A3(new_n860), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT111), .B1(new_n685), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n685), .A2(KEYINPUT111), .A3(new_n874), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n866), .A2(new_n872), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n847), .B1(new_n856), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n762), .A2(new_n637), .A3(new_n752), .A4(new_n753), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n771), .B1(new_n881), .B2(new_n707), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n646), .A2(new_n637), .A3(new_n752), .A4(new_n753), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n707), .A2(new_n883), .A3(new_n388), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n627), .A2(KEYINPUT110), .A3(new_n861), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT110), .B1(new_n627), .B2(new_n861), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n885), .B(new_n760), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n685), .A2(KEYINPUT111), .A3(new_n874), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n875), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n794), .A2(new_n797), .A3(new_n801), .A4(new_n871), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT113), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n855), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n775), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n708), .B2(new_n718), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT113), .B1(new_n897), .B2(new_n852), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n894), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(new_n899), .A3(KEYINPUT53), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n880), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n856), .A2(new_n879), .A3(new_n847), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n906), .B2(new_n847), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n907), .B2(new_n901), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n805), .A2(new_n618), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n759), .A2(new_n770), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n636), .A4(new_n722), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT50), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n759), .A2(new_n619), .A3(new_n808), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n388), .A3(new_n732), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n734), .A2(new_n740), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n805), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n914), .A2(new_n915), .B1(new_n916), .B2(new_n774), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n749), .A2(new_n492), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n835), .B1(new_n709), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n770), .A3(new_n808), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n912), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n909), .A2(new_n754), .A3(new_n770), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n616), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n785), .A2(new_n389), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n916), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT48), .Z(new_n930));
  AOI211_X1 g744(.A(new_n927), .B(new_n930), .C1(new_n859), .C2(new_n914), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n924), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n908), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  INV_X1    g747(.A(new_n732), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n918), .B(KEYINPUT49), .Z(new_n935));
  NOR4_X1   g749(.A1(new_n804), .A2(new_n388), .A3(new_n636), .A4(new_n709), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n722), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT109), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n933), .A2(new_n938), .ZN(G75));
  AOI21_X1  g753(.A(new_n297), .B1(new_n880), .B2(new_n900), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(new_n450), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n426), .A2(new_n434), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT114), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n432), .B(KEYINPUT55), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n941), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n321), .A2(G952), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT115), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(G51));
  AND2_X1   g764(.A1(new_n940), .A2(new_n818), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n902), .A2(KEYINPUT116), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n880), .A2(new_n900), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT116), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n880), .A2(new_n900), .A3(new_n955), .A4(new_n901), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n499), .B(KEYINPUT57), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n748), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n951), .B1(new_n959), .B2(KEYINPUT117), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT117), .ZN(new_n961));
  INV_X1    g775(.A(new_n958), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n901), .B1(new_n880), .B2(new_n900), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n880), .A2(new_n900), .A3(new_n901), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n955), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n965), .B2(new_n952), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n961), .B1(new_n966), .B2(new_n748), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n947), .B1(new_n960), .B2(new_n967), .ZN(G54));
  NAND3_X1  g782(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(new_n660), .ZN(new_n970));
  INV_X1    g784(.A(new_n947), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n660), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT118), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n970), .A2(KEYINPUT118), .A3(new_n971), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G60));
  AND2_X1   g791(.A1(new_n639), .A2(new_n641), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n644), .B(KEYINPUT59), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n908), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n957), .A2(new_n979), .A3(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n949), .ZN(G63));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT60), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n953), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n949), .B1(new_n986), .B2(new_n690), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n676), .A2(new_n677), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n953), .A2(new_n988), .A3(new_n985), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT119), .ZN(new_n990));
  AOI22_X1  g804(.A1(new_n987), .A2(new_n989), .B1(new_n990), .B2(KEYINPUT61), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G66));
  OAI21_X1  g807(.A(G953), .B1(new_n622), .B2(new_n430), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n888), .A2(new_n890), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n943), .B1(G898), .B2(new_n321), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G69));
  OAI21_X1  g812(.A(new_n281), .B1(KEYINPUT30), .B2(new_n252), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n547), .B1(new_n338), .B2(new_n548), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT120), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n897), .A2(new_n743), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(KEYINPUT62), .A3(new_n738), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g821(.A(new_n738), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n859), .A2(new_n873), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1011), .A2(new_n724), .A3(new_n869), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n318), .A3(new_n389), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT121), .B1(new_n828), .B2(new_n1013), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n828), .A2(KEYINPUT121), .A3(new_n1013), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1010), .B(new_n845), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1003), .B1(new_n1016), .B2(new_n321), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT122), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n828), .A2(new_n1005), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1018), .B1(new_n828), .B2(new_n1005), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n850), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n823), .A2(new_n827), .A3(new_n1023), .A4(new_n928), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1024), .A2(new_n798), .A3(new_n801), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n845), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT123), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1021), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1019), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1024), .A2(new_n798), .A3(new_n801), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1030), .B1(new_n842), .B2(new_n844), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT123), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1027), .A2(new_n321), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1001), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1035), .B1(G900), .B2(G953), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1017), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n1037), .A2(KEYINPUT124), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1038), .A2(KEYINPUT124), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1038), .A2(KEYINPUT124), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1039), .A2(new_n1042), .ZN(G72));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1044), .B(KEYINPUT126), .ZN(new_n1045));
  XNOR2_X1  g859(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1046));
  XNOR2_X1  g860(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT127), .Z(new_n1048));
  INV_X1    g862(.A(new_n995), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1048), .B1(new_n1016), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1050), .A2(new_n278), .A3(new_n726), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n271), .A2(new_n279), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1047), .B1(new_n306), .B2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g867(.A(new_n1051), .B(new_n971), .C1(new_n907), .C2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1027), .A2(new_n995), .A3(new_n1033), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1055), .A2(new_n1048), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n726), .A2(new_n278), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(G57));
endmodule


