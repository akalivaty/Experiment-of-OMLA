//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR3_X1   g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n210), .A2(new_n214), .A3(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(KEYINPUT76), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n248), .A2(new_n252), .B1(new_n251), .B2(new_n245), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT74), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G58), .A2(G68), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT73), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT73), .B1(G58), .B2(G68), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n257), .A2(new_n201), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n259), .B2(new_n212), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n255), .B(new_n256), .ZN(new_n261));
  OAI211_X1 g0061(.A(KEYINPUT74), .B(G20), .C1(new_n261), .C2(new_n201), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G159), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G68), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n263), .A2(new_n265), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT16), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n250), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n263), .A2(new_n276), .A3(KEYINPUT16), .A4(new_n265), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n253), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n267), .A2(G226), .A3(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n267), .A2(G223), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G87), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT68), .A2(G41), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT68), .A2(G41), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  AND2_X1   g0098(.A1(G1), .A2(G13), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n287), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n288), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n297), .A2(new_n300), .B1(new_n302), .B2(G232), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n290), .A2(new_n291), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT75), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n290), .A2(new_n303), .A3(KEYINPUT75), .A4(new_n291), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n290), .A2(new_n303), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT18), .B1(new_n281), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n277), .A2(new_n278), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n249), .A2(new_n213), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n280), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n253), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT18), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n306), .A2(new_n307), .B1(new_n310), .B2(new_n309), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n243), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n281), .B2(new_n312), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n309), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n290), .B2(new_n303), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n316), .A2(new_n329), .A3(new_n317), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n281), .A2(KEYINPUT17), .A3(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n324), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n322), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n273), .A2(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G222), .ZN(new_n337));
  INV_X1    g0137(.A(G77), .ZN(new_n338));
  INV_X1    g0138(.A(G223), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n267), .A2(G1698), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n337), .B1(new_n338), .B2(new_n267), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n289), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n297), .A2(new_n300), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(G226), .B2(new_n302), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n310), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n212), .A2(G33), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n245), .A2(new_n349), .B1(G150), .B2(new_n264), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n203), .A2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n315), .ZN(new_n353));
  INV_X1    g0153(.A(new_n251), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n315), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(G50), .A3(new_n247), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n353), .B(new_n356), .C1(G50), .C2(new_n251), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n347), .B(new_n357), .C1(G179), .C2(new_n346), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n342), .A2(new_n345), .A3(G190), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT70), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT10), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n357), .A2(KEYINPUT9), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(KEYINPUT9), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n362), .A2(new_n363), .B1(G200), .B2(new_n346), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(new_n364), .B2(new_n360), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n358), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n355), .A2(G68), .A3(new_n247), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n368), .B(KEYINPUT72), .Z(new_n369));
  AOI22_X1  g0169(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n338), .B2(new_n348), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(new_n315), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n354), .A2(new_n216), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n376));
  AND4_X1   g0176(.A1(new_n369), .A2(new_n373), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT71), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n336), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n289), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n302), .A2(G238), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n343), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n288), .B1(new_n380), .B2(new_n381), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT13), .B1(new_n389), .B2(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(G169), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(G179), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n391), .B2(G169), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n378), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n377), .B1(new_n391), .B2(new_n325), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n327), .B1(new_n388), .B2(new_n390), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n245), .A2(new_n264), .B1(G20), .B2(G77), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n349), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n250), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n355), .A2(G77), .A3(new_n247), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G77), .B2(new_n251), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n302), .A2(G244), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n336), .A2(G232), .ZN(new_n413));
  INV_X1    g0213(.A(G107), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n414), .B2(new_n267), .C1(new_n215), .C2(new_n340), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n344), .B(new_n412), .C1(new_n415), .C2(new_n289), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(G169), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT69), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n291), .ZN(new_n420));
  OAI211_X1 g0220(.A(KEYINPUT69), .B(new_n411), .C1(new_n416), .C2(G169), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(G190), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n410), .C1(new_n327), .C2(new_n416), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OR4_X1    g0225(.A1(new_n335), .A2(new_n367), .A3(new_n402), .A4(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT77), .B1(new_n273), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G283), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT77), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n267), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n270), .A2(new_n272), .A3(G250), .A4(G1698), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n428), .A2(new_n429), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n270), .A2(new_n272), .A3(G244), .A4(new_n283), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT4), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n289), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(KEYINPUT68), .A2(G41), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT5), .B1(new_n440), .B2(new_n292), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT5), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n246), .B(G45), .C1(new_n442), .C2(G41), .ZN(new_n443));
  OAI211_X1 g0243(.A(G257), .B(new_n288), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n293), .B2(new_n294), .ZN(new_n445));
  INV_X1    g0245(.A(new_n443), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n300), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n439), .A2(new_n291), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n439), .A2(KEYINPUT79), .A3(new_n291), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT78), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n433), .A2(new_n429), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(new_n437), .A3(new_n428), .A4(new_n432), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n455), .B(new_n448), .C1(new_n289), .C2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT78), .B1(new_n439), .B2(new_n449), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n310), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n414), .A2(KEYINPUT6), .A3(G97), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n414), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G97), .A2(G107), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(KEYINPUT6), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n264), .A2(G77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n414), .B1(new_n268), .B2(new_n274), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n315), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n354), .A2(new_n462), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n250), .B(new_n251), .C1(G1), .C2(new_n269), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n454), .A2(new_n460), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n439), .A2(new_n449), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n455), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n439), .A2(KEYINPUT78), .A3(new_n449), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(G190), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(G200), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n270), .A2(new_n272), .A3(G264), .A4(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n270), .A2(new_n272), .A3(G257), .A4(new_n283), .ZN(new_n489));
  INV_X1    g0289(.A(G303), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(new_n267), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(new_n289), .ZN(new_n492));
  OAI211_X1 g0292(.A(G270), .B(new_n288), .C1(new_n441), .C2(new_n443), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n447), .ZN(new_n494));
  OAI21_X1  g0294(.A(G169), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n354), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n473), .B2(new_n496), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n249), .A2(new_n213), .B1(G20), .B2(new_n496), .ZN(new_n499));
  AOI21_X1  g0299(.A(G20), .B1(G33), .B2(G283), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n269), .A2(G97), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT81), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT81), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT20), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n487), .B1(new_n495), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT82), .B(new_n487), .C1(new_n495), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n491), .A2(new_n289), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(G179), .A3(new_n447), .A4(new_n493), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n495), .B2(new_n487), .ZN(new_n516));
  INV_X1    g0316(.A(new_n508), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n447), .A3(new_n493), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G200), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n508), .C1(new_n325), .C2(new_n519), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G264), .B(new_n288), .C1(new_n441), .C2(new_n443), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n445), .A2(new_n446), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT85), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(G264), .A4(new_n288), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n267), .A2(G250), .A3(new_n283), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n525), .A2(new_n528), .B1(new_n289), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(G179), .A3(new_n447), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n528), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n289), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(new_n447), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n534), .B(new_n535), .C1(new_n538), .C2(new_n310), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(KEYINPUT86), .A3(G179), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT25), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n251), .B2(G107), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n251), .A2(new_n541), .A3(G107), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n473), .A2(new_n414), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n270), .A2(new_n272), .A3(new_n212), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n267), .A2(new_n547), .A3(new_n212), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G116), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(G20), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n212), .B2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n414), .A2(KEYINPUT23), .A3(G20), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT84), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT84), .A4(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(KEYINPUT24), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n315), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n546), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n539), .A2(new_n540), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n533), .A2(new_n325), .A3(new_n447), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n538), .B2(G200), .ZN(new_n570));
  INV_X1    g0370(.A(new_n566), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n545), .B1(new_n571), .B2(new_n562), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n212), .ZN(new_n576));
  INV_X1    g0376(.A(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n464), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n270), .A2(new_n272), .A3(new_n212), .A4(G68), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n348), .B2(new_n462), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n315), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n404), .A2(new_n354), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G250), .B1(new_n296), .B2(G1), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n299), .B2(new_n287), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT80), .ZN(new_n589));
  AND2_X1   g0389(.A1(G33), .A2(G41), .ZN(new_n590));
  OAI21_X1  g0390(.A(G274), .B1(new_n590), .B2(new_n213), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n246), .A2(G45), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n296), .A2(G1), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n300), .A2(KEYINPUT80), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n270), .A2(new_n272), .A3(G244), .A4(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n270), .A2(new_n272), .A3(G238), .A4(new_n283), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n552), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n289), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(G190), .A3(new_n600), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n473), .A2(new_n577), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n586), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n596), .A2(new_n291), .A3(new_n600), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n355), .B(new_n405), .C1(G1), .C2(new_n269), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n584), .A2(new_n607), .A3(new_n585), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n310), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n603), .A2(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n486), .A2(new_n523), .A3(new_n574), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n426), .A2(new_n612), .ZN(G372));
  NAND2_X1  g0413(.A1(new_n332), .A2(new_n333), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n614), .B(new_n400), .C1(new_n397), .C2(new_n422), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n313), .A2(new_n321), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n366), .B2(new_n365), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n358), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n593), .A2(new_n595), .ZN(new_n620));
  INV_X1    g0420(.A(new_n588), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT87), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT87), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n623), .B(new_n588), .C1(new_n593), .C2(new_n595), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n600), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n310), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT88), .B1(new_n626), .B2(new_n606), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n596), .A2(new_n291), .A3(new_n600), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n625), .C2(new_n310), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n608), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(G200), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n570), .A2(new_n572), .B1(new_n603), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n634), .A2(new_n477), .A3(new_n484), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n568), .A2(new_n518), .A3(new_n513), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n603), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n600), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT80), .B1(new_n300), .B2(new_n594), .ZN(new_n641));
  AND4_X1   g0441(.A1(KEYINPUT80), .A2(new_n288), .A3(G274), .A4(new_n594), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n621), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n623), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n596), .A2(KEYINPUT87), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n606), .B1(new_n646), .B2(G169), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n628), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n626), .A2(KEYINPUT88), .A3(new_n606), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n650), .B2(new_n608), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n454), .A2(new_n460), .A3(new_n476), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT26), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n611), .A2(new_n454), .A3(new_n460), .A4(new_n476), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n637), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n619), .B1(new_n426), .B2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n246), .A2(new_n212), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n508), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n522), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n513), .A2(new_n518), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n667), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT89), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(G330), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n574), .B1(new_n572), .B2(new_n666), .ZN(new_n677));
  INV_X1    g0477(.A(new_n568), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n665), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n665), .B1(new_n513), .B2(new_n518), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n574), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n568), .B2(new_n665), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n681), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n208), .ZN(new_n687));
  INV_X1    g0487(.A(new_n295), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n578), .A2(G116), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n246), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n211), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n689), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  NAND3_X1  g0495(.A1(new_n631), .A2(new_n652), .A3(new_n638), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n656), .B1(new_n696), .B2(new_n655), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n568), .A2(new_n518), .A3(new_n513), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n634), .A2(new_n477), .A3(new_n484), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n631), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n666), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(KEYINPUT26), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n632), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n477), .A2(new_n484), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n636), .A2(new_n573), .A3(new_n631), .A4(new_n638), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n704), .B(new_n706), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT94), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n703), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n712), .A2(KEYINPUT94), .A3(KEYINPUT29), .A4(new_n666), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n666), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n536), .A2(new_n537), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n720), .A2(new_n604), .A3(new_n515), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n479), .A3(new_n480), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n538), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n519), .A2(new_n291), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n478), .A3(new_n625), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT90), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT30), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n721), .A2(KEYINPUT90), .A3(new_n479), .A4(new_n480), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n724), .B1(new_n732), .B2(KEYINPUT91), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n479), .A2(new_n480), .ZN(new_n734));
  INV_X1    g0534(.A(new_n515), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n533), .A3(new_n600), .A4(new_n596), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n729), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n723), .A3(new_n731), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(KEYINPUT91), .A3(new_n727), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n719), .B1(new_n733), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(new_n727), .A3(new_n724), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT92), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n738), .A2(new_n724), .A3(KEYINPUT92), .A4(new_n727), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n666), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n568), .A2(new_n573), .A3(new_n611), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n746), .A2(new_n485), .A3(new_n522), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n718), .B1(new_n747), .B2(new_n666), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n740), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n717), .B1(G330), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n695), .B1(new_n750), .B2(G1), .ZN(G364));
  NAND2_X1  g0551(.A1(new_n672), .A2(new_n674), .ZN(new_n752));
  INV_X1    g0552(.A(G330), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n689), .ZN(new_n755));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n246), .B1(new_n757), .B2(G45), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n675), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n213), .B1(G20), .B2(new_n310), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n212), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n325), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n414), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n212), .A2(new_n291), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n766), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n325), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G58), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n267), .B1(new_n338), .B2(new_n768), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n325), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n212), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n765), .B(new_n773), .C1(G97), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n763), .A2(new_n767), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT32), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n778), .A2(KEYINPUT32), .A3(new_n779), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(G87), .B2(new_n783), .ZN(new_n784));
  AND3_X1   g0584(.A1(new_n777), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT98), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n769), .B2(new_n327), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n766), .A2(KEYINPUT98), .A3(G200), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(G190), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n787), .A2(new_n325), .A3(new_n788), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n785), .B1(new_n202), .B2(new_n793), .C1(new_n216), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n775), .A2(new_n796), .B1(new_n782), .B2(new_n490), .ZN(new_n797));
  INV_X1    g0597(.A(new_n778), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n267), .B1(new_n798), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n768), .C1(new_n771), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n764), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n797), .B(new_n802), .C1(G283), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(G326), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n805), .C1(new_n794), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n762), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n761), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n241), .A2(G45), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n687), .A2(new_n267), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n296), .B2(new_n693), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n687), .A2(new_n273), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(G355), .B(KEYINPUT95), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n821), .B1(G116), .B2(new_n208), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT96), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n815), .A2(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n814), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n809), .A2(new_n826), .A3(new_n759), .ZN(new_n827));
  INV_X1    g0627(.A(new_n812), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n671), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n760), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n411), .A2(new_n665), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n422), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n422), .A2(new_n424), .A3(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n810), .ZN(new_n837));
  INV_X1    g0637(.A(new_n759), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n761), .A2(new_n810), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(G77), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n776), .A2(G97), .B1(new_n803), .B2(G87), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n414), .B2(new_n782), .ZN(new_n843));
  INV_X1    g0643(.A(new_n768), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n267), .B1(new_n844), .B2(G116), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n800), .B2(new_n778), .C1(new_n771), .C2(new_n796), .ZN(new_n846));
  INV_X1    g0646(.A(new_n794), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n843), .B(new_n846), .C1(G283), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n490), .B2(new_n793), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n764), .A2(new_n216), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n273), .B(new_n850), .C1(G132), .C2(new_n798), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n776), .A2(G58), .B1(new_n783), .B2(G50), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n770), .A2(G143), .B1(G159), .B2(new_n844), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n794), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n792), .B2(G137), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n851), .B(new_n852), .C1(new_n856), .C2(KEYINPUT34), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n841), .B1(new_n859), .B2(new_n761), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n837), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n835), .B(KEYINPUT101), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n701), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n425), .A2(new_n665), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT102), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(new_n697), .C2(new_n700), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n865), .B1(new_n657), .B2(new_n864), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n749), .A2(G330), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n759), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n870), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n861), .B1(new_n873), .B2(new_n875), .ZN(G384));
  NOR2_X1   g0676(.A1(new_n757), .A2(new_n246), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n426), .B1(new_n715), .B2(new_n716), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n618), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT107), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n422), .A2(new_n665), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n868), .B2(new_n867), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n281), .A2(new_n663), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n322), .B2(new_n334), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n330), .B1(new_n281), .B2(new_n312), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n886), .B2(new_n884), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n318), .A2(new_n320), .ZN(new_n888));
  INV_X1    g0688(.A(new_n663), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n318), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n888), .A2(new_n890), .A3(new_n330), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n885), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n378), .A2(new_n665), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n397), .B2(new_n401), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n397), .A2(new_n401), .A3(new_n899), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n883), .A2(new_n898), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n616), .A2(new_n663), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n885), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(new_n891), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n886), .B2(new_n884), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n892), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n884), .B1(new_n616), .B2(new_n614), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n906), .B1(new_n913), .B2(KEYINPUT39), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n397), .A2(new_n665), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n905), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n904), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n880), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT92), .B1(new_n732), .B2(new_n724), .ZN(new_n919));
  INV_X1    g0719(.A(new_n744), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n665), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT31), .B1(new_n612), .B2(new_n665), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n743), .A2(new_n744), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n925), .B2(new_n719), .ZN(new_n926));
  INV_X1    g0726(.A(new_n719), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT108), .B(new_n927), .C1(new_n743), .C2(new_n744), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n923), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n836), .B1(new_n902), .B2(new_n901), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n898), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n912), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n934), .B2(new_n897), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n719), .B1(new_n919), .B2(new_n920), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT108), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n925), .A2(new_n924), .A3(new_n719), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n426), .B1(new_n923), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n753), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n937), .B2(new_n942), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n877), .B1(new_n918), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n918), .B2(new_n944), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n213), .A2(new_n212), .A3(new_n496), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n466), .B(KEYINPUT104), .Z(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT35), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  NOR3_X1   g0753(.A1(new_n261), .A2(new_n338), .A3(new_n211), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n954), .A2(new_n955), .B1(new_n202), .B2(G68), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(G1), .A3(new_n756), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n946), .A2(new_n953), .A3(new_n958), .ZN(G367));
  OAI211_X1 g0759(.A(new_n707), .B(new_n709), .C1(new_n482), .C2(new_n666), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n477), .A2(new_n666), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n683), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n477), .B1(new_n960), .B2(new_n568), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n965), .A2(KEYINPUT42), .B1(new_n967), .B2(new_n666), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n666), .B1(new_n586), .B2(new_n602), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n632), .A2(new_n639), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n632), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n966), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n963), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n681), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n689), .B(KEYINPUT41), .Z(new_n981));
  INV_X1    g0781(.A(new_n717), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n680), .A2(new_n682), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n964), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n675), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n870), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT111), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n750), .A2(KEYINPUT111), .A3(new_n985), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n684), .A2(new_n960), .A3(new_n962), .ZN(new_n990));
  NOR2_X1   g0790(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n978), .B2(new_n684), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n963), .A2(new_n685), .A3(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n999), .A3(new_n681), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n995), .A2(new_n999), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n681), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(KEYINPUT110), .A3(new_n1003), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n988), .A2(new_n989), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n981), .B1(new_n1007), .B2(new_n750), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n758), .B(KEYINPUT112), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n980), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n814), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n208), .B2(new_n404), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n817), .A2(new_n233), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n838), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n776), .A2(G68), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n772), .B2(new_n782), .C1(new_n338), .C2(new_n764), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n273), .B1(new_n844), .B2(G50), .ZN(new_n1017));
  INV_X1    g0817(.A(G137), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n778), .C1(new_n771), .C2(new_n854), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(G159), .C2(new_n847), .ZN(new_n1020));
  INV_X1    g0820(.A(G143), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n793), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n782), .A2(new_n496), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT46), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n764), .A2(new_n462), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G107), .B2(new_n776), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n798), .A2(G317), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n267), .B1(new_n844), .B2(G283), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1024), .B(new_n1029), .C1(G294), .C2(new_n847), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n792), .A2(G311), .B1(G303), .B2(new_n770), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(new_n1031), .B2(KEYINPUT113), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(KEYINPUT113), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1022), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1014), .B1(new_n1035), .B2(new_n761), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n970), .A2(new_n812), .A3(new_n971), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1010), .A2(new_n1038), .ZN(G387));
  AND2_X1   g0839(.A1(new_n989), .A2(new_n988), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n689), .B1(new_n750), .B2(new_n985), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n985), .A2(new_n1009), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n244), .A2(G50), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT50), .Z(new_n1046));
  OAI211_X1 g0846(.A(new_n690), .B(new_n296), .C1(new_n216), .C2(new_n338), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n816), .B1(new_n1046), .B2(new_n1047), .C1(new_n230), .C2(new_n296), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n819), .A2(new_n691), .B1(new_n414), .B2(new_n687), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(KEYINPUT114), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(KEYINPUT114), .B2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n838), .B1(new_n1051), .B2(new_n814), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G68), .A2(new_n844), .B1(new_n798), .B2(G150), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n267), .C1(new_n202), .C2(new_n771), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n775), .A2(new_n404), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n782), .A2(new_n338), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1054), .A2(new_n1025), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n244), .B2(new_n794), .C1(new_n779), .C2(new_n793), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n267), .B1(new_n798), .B2(G326), .ZN(new_n1059));
  INV_X1    g0859(.A(G283), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n775), .A2(new_n1060), .B1(new_n782), .B2(new_n796), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n770), .A2(G317), .B1(G303), .B2(new_n844), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n800), .B2(new_n794), .C1(new_n793), .C2(new_n801), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1059), .B1(new_n496), .B2(new_n764), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1052), .B1(new_n1070), .B2(new_n761), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n680), .B2(new_n828), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1044), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1043), .A2(new_n1074), .ZN(G393));
  AND2_X1   g0875(.A1(new_n1004), .A2(new_n1000), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1007), .B(new_n689), .C1(new_n1040), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1009), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n792), .A2(G150), .B1(G159), .B2(new_n770), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n794), .A2(new_n202), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n267), .B1(new_n778), .B2(new_n1021), .C1(new_n244), .C2(new_n768), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n775), .A2(new_n338), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n216), .B2(new_n782), .C1(new_n577), .C2(new_n764), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n792), .A2(G317), .B1(G311), .B2(new_n770), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n794), .A2(new_n490), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n273), .B1(new_n778), .B2(new_n801), .C1(new_n796), .C2(new_n768), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n765), .B1(G283), .B2(new_n783), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n496), .B2(new_n775), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n761), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n238), .A2(new_n817), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n814), .B1(G97), .B2(new_n687), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n759), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1095), .B(new_n1099), .C1(new_n963), .C2(new_n828), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1077), .A2(new_n1078), .A3(new_n1100), .ZN(G390));
  OAI21_X1  g0901(.A(new_n915), .B1(new_n907), .B2(new_n912), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n712), .A2(new_n666), .A3(new_n835), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n882), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n903), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n749), .A2(G330), .A3(new_n835), .A4(new_n903), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n864), .B1(new_n697), .B2(new_n700), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT102), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n881), .B1(new_n1109), .B2(new_n866), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n903), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n915), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1105), .B(new_n1107), .C1(new_n914), .C2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n929), .A2(G330), .A3(new_n930), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n914), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1105), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n335), .A2(new_n367), .A3(new_n402), .A4(new_n425), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n929), .A2(G330), .A3(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n619), .B(new_n1120), .C1(new_n982), .C2(new_n426), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n862), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n929), .A3(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1111), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1104), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n1106), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1111), .B1(new_n870), .B2(new_n836), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1114), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n883), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1121), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n755), .B1(new_n1118), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n915), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n883), .B2(new_n903), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n914), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1106), .B(new_n1116), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1105), .B1(new_n1112), .B2(new_n914), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n1114), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n929), .A2(G330), .A3(new_n1119), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1138), .A2(new_n878), .A3(new_n618), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1106), .A2(new_n1125), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1111), .B2(new_n1123), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1110), .B1(new_n1127), .B2(new_n1114), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1137), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1131), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1134), .A2(new_n811), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n771), .A2(new_n496), .B1(new_n768), .B2(new_n462), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n267), .B(new_n1149), .C1(G294), .C2(new_n798), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n850), .B(new_n1083), .C1(G87), .C2(new_n783), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n414), .C2(new_n794), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G283), .B2(new_n792), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n847), .A2(G137), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n782), .A2(new_n854), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n776), .A2(G159), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n770), .A2(G132), .B1(new_n844), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n273), .B1(new_n798), .B2(G125), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n202), .B2(new_n764), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT118), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1161), .B(new_n1164), .C1(G128), .C2(new_n792), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n761), .B1(new_n1153), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n838), .C1(new_n245), .C2(new_n840), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1148), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1135), .B(new_n1009), .C1(new_n1114), .C2(new_n1136), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT117), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1114), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(KEYINPUT117), .A3(new_n1009), .A4(new_n1135), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1168), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1147), .A2(new_n1176), .ZN(G378));
  OAI21_X1  g0977(.A(new_n838), .B1(G50), .B2(new_n840), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n295), .B2(new_n273), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n803), .A2(G58), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1015), .B(new_n1181), .C1(new_n338), .C2(new_n782), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n771), .A2(new_n414), .B1(new_n778), .B2(new_n1060), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n295), .B(new_n273), .C1(new_n768), .C2(new_n404), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n462), .B2(new_n794), .C1(new_n793), .C2(new_n496), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G132), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n794), .A2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n770), .A2(G128), .B1(G137), .B2(new_n844), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n854), .B2(new_n775), .C1(new_n782), .C2(new_n1158), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G125), .C2(new_n792), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n779), .B2(new_n764), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT119), .Z(new_n1198));
  INV_X1    g0998(.A(KEYINPUT59), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .C1(new_n1195), .C2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1178), .B1(new_n1201), .B2(new_n761), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n357), .A2(new_n889), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n367), .B(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1204), .B(new_n1205), .Z(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1202), .B1(new_n1207), .B2(new_n811), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT120), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n903), .A2(new_n835), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n941), .B2(new_n923), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT40), .B1(new_n1211), .B2(new_n898), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n936), .A2(G330), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n933), .A2(new_n1206), .A3(G330), .A4(new_n936), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(KEYINPUT121), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n917), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n917), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1218), .A2(new_n1214), .A3(KEYINPUT121), .A4(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1209), .B1(new_n1220), .B2(new_n1009), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1218), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1214), .A2(new_n917), .A3(new_n1215), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT57), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1121), .B1(new_n1118), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n689), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1139), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1221), .B1(new_n1228), .B2(new_n1230), .ZN(G375));
  NAND2_X1  g1031(.A1(new_n1111), .A2(new_n810), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1181), .B1(new_n779), .B2(new_n782), .C1(new_n202), .C2(new_n775), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n273), .B1(new_n798), .B2(G128), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n854), .B2(new_n768), .C1(new_n771), .C2(new_n1018), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(new_n847), .C2(new_n1159), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1189), .B2(new_n793), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n775), .A2(new_n404), .B1(new_n782), .B2(new_n462), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G107), .A2(new_n844), .B1(new_n798), .B2(G303), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1060), .B2(new_n771), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G116), .C2(new_n847), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n273), .B1(new_n764), .B2(new_n338), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT122), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(new_n796), .C2(new_n793), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n762), .B1(new_n1237), .B2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n759), .B(new_n1245), .C1(new_n216), .C2(new_n839), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT123), .Z(new_n1247));
  AOI22_X1  g1047(.A1(new_n1226), .A2(new_n1009), .B1(new_n1232), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1126), .A2(new_n1121), .A3(new_n1129), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n981), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1143), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G381));
  NAND3_X1  g1052(.A1(new_n1043), .A2(new_n830), .A3(new_n1074), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G384), .ZN(new_n1254));
  AOI211_X1 g1054(.A(G390), .B(G381), .C1(new_n1254), .C2(KEYINPUT124), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G387), .A2(G378), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(KEYINPUT124), .C2(new_n1254), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(G375), .ZN(G407));
  OAI21_X1  g1058(.A(new_n689), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT116), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1137), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1168), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n664), .A2(G213), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT125), .Z(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G375), .C2(new_n1270), .ZN(G409));
  AND2_X1   g1071(.A1(new_n1010), .A2(new_n1038), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT127), .B1(new_n1272), .B2(G390), .ZN(new_n1273));
  OAI21_X1  g1073(.A(G396), .B1(new_n1042), .B2(new_n1073), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1253), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(G390), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G390), .B1(new_n1010), .B2(new_n1038), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1273), .A2(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G390), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G387), .A2(new_n1281), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(new_n1282), .A2(new_n1278), .A3(KEYINPUT127), .A4(new_n1275), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1221), .C1(new_n1230), .C2(new_n1228), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1214), .A2(new_n917), .A3(new_n1215), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n917), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1209), .B1(new_n1289), .B2(new_n1009), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1220), .A2(new_n1250), .A3(new_n1229), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1267), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1286), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1269), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  XOR2_X1   g1096(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n1297));
  NAND2_X1  g1097(.A1(new_n1249), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1126), .A2(new_n1121), .A3(new_n1129), .A4(KEYINPUT60), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n689), .A3(new_n1143), .A4(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(G384), .A3(new_n1248), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G384), .B1(new_n1300), .B2(new_n1248), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1285), .B1(new_n1296), .B2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G2897), .B(new_n1269), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1303), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1269), .A2(G2897), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1301), .A3(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1269), .B1(new_n1286), .B2(new_n1293), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1304), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1284), .A2(new_n1306), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1313), .A2(new_n1316), .A3(new_n1304), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1313), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(new_n1313), .B2(new_n1304), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1317), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1322), .B2(new_n1284), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1267), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1286), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1280), .A2(new_n1283), .A3(new_n1304), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1278), .A2(new_n1327), .ZN(new_n1328));
  OAI22_X1  g1128(.A1(new_n1328), .A2(new_n1275), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1277), .A2(new_n1279), .A3(new_n1327), .A4(new_n1276), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1305), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1325), .B1(new_n1326), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1304), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1330), .A3(new_n1305), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1333), .A2(new_n1286), .A3(new_n1324), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1332), .A2(new_n1335), .ZN(G402));
endmodule


