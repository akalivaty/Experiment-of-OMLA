

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582;

  NAND2_X1 U319 ( .A1(n472), .A2(n471), .ZN(n486) );
  NOR2_X1 U320 ( .A1(n580), .A2(n487), .ZN(n489) );
  XOR2_X1 U321 ( .A(n349), .B(n348), .Z(n287) );
  XOR2_X1 U322 ( .A(G127GAT), .B(KEYINPUT81), .Z(n288) );
  XOR2_X1 U323 ( .A(n415), .B(n315), .Z(n289) );
  INV_X1 U324 ( .A(KEYINPUT99), .ZN(n469) );
  XNOR2_X1 U325 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U326 ( .A(n350), .B(n287), .ZN(n351) );
  XNOR2_X1 U327 ( .A(n316), .B(n289), .ZN(n317) );
  XNOR2_X1 U328 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U329 ( .A(n447), .B(KEYINPUT119), .ZN(n448) );
  NOR2_X1 U330 ( .A1(n464), .A2(n528), .ZN(n461) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U332 ( .A(KEYINPUT38), .B(n491), .Z(n497) );
  XNOR2_X1 U333 ( .A(n453), .B(KEYINPUT122), .ZN(n454) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  XOR2_X1 U336 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XNOR2_X1 U337 ( .A(n441), .B(n396), .ZN(n291) );
  AND2_X1 U338 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U340 ( .A(KEYINPUT10), .B(KEYINPUT78), .Z(n293) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G106GAT), .ZN(n292) );
  XOR2_X1 U342 ( .A(n293), .B(n292), .Z(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n300) );
  XOR2_X1 U344 ( .A(G43GAT), .B(G134GAT), .Z(n318) );
  XOR2_X1 U345 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n297) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n318), .B(n298), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n301), .B(G92GAT), .Z(n305) );
  XOR2_X1 U351 ( .A(G29GAT), .B(KEYINPUT7), .Z(n303) );
  XNOR2_X1 U352 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n336) );
  XNOR2_X1 U354 ( .A(n336), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n552) );
  INV_X1 U356 ( .A(n552), .ZN(n536) );
  XOR2_X1 U357 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U358 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U360 ( .A(n308), .B(G183GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G176GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n390) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G71GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n311), .B(G120GAT), .ZN(n347) );
  XNOR2_X1 U365 ( .A(G15GAT), .B(n347), .ZN(n316) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n288), .B(n312), .ZN(n415) );
  XOR2_X1 U368 ( .A(KEYINPUT20), .B(KEYINPUT66), .Z(n314) );
  NAND2_X1 U369 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(n317), .B(KEYINPUT83), .Z(n320) );
  XNOR2_X1 U372 ( .A(n318), .B(G190GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X2 U374 ( .A(n390), .B(n321), .Z(n519) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n323) );
  XNOR2_X1 U376 ( .A(KEYINPUT68), .B(KEYINPUT73), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n330) );
  XOR2_X1 U378 ( .A(G197GAT), .B(G36GAT), .Z(n325) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(G43GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U381 ( .A(n326), .B(G113GAT), .Z(n328) );
  XOR2_X1 U382 ( .A(G141GAT), .B(G22GAT), .Z(n442) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(n442), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n340) );
  XOR2_X1 U386 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n332) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U389 ( .A(n333), .B(KEYINPUT30), .Z(n338) );
  XOR2_X1 U390 ( .A(G1GAT), .B(G8GAT), .Z(n335) );
  XNOR2_X1 U391 ( .A(G15GAT), .B(KEYINPUT72), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n369) );
  XNOR2_X1 U393 ( .A(n336), .B(n369), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n568) );
  XOR2_X1 U396 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n342) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n354) );
  XNOR2_X1 U399 ( .A(G204GAT), .B(G92GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n343), .B(G64GAT), .ZN(n389) );
  XOR2_X1 U401 ( .A(G85GAT), .B(G57GAT), .Z(n416) );
  XOR2_X1 U402 ( .A(n389), .B(n416), .Z(n345) );
  NAND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n352) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n346), .B(G148GAT), .ZN(n436) );
  XNOR2_X1 U407 ( .A(n347), .B(n436), .ZN(n350) );
  XOR2_X1 U408 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n349) );
  XNOR2_X1 U409 ( .A(KEYINPUT13), .B(KEYINPUT76), .ZN(n348) );
  XOR2_X1 U410 ( .A(n354), .B(n353), .Z(n573) );
  XOR2_X1 U411 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n355) );
  XNOR2_X1 U412 ( .A(n573), .B(n355), .ZN(n499) );
  NOR2_X1 U413 ( .A1(n568), .A2(n499), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n356), .B(KEYINPUT46), .ZN(n374) );
  XOR2_X1 U415 ( .A(G64GAT), .B(G127GAT), .Z(n358) );
  XNOR2_X1 U416 ( .A(G183GAT), .B(G71GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n360) );
  XNOR2_X1 U419 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n373) );
  XOR2_X1 U422 ( .A(G211GAT), .B(G155GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(G22GAT), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U425 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n366) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(n368), .B(n367), .Z(n371) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT14), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n562) );
  NOR2_X1 U432 ( .A1(n374), .A2(n562), .ZN(n375) );
  NAND2_X1 U433 ( .A1(n375), .A2(n552), .ZN(n378) );
  INV_X1 U434 ( .A(n378), .ZN(n377) );
  XOR2_X1 U435 ( .A(KEYINPUT111), .B(KEYINPUT47), .Z(n379) );
  INV_X1 U436 ( .A(n379), .ZN(n376) );
  NAND2_X1 U437 ( .A1(n377), .A2(n376), .ZN(n381) );
  NAND2_X1 U438 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U439 ( .A1(n381), .A2(n380), .ZN(n387) );
  INV_X1 U440 ( .A(n568), .ZN(n555) );
  XNOR2_X1 U441 ( .A(n552), .B(KEYINPUT36), .ZN(n580) );
  INV_X1 U442 ( .A(n562), .ZN(n577) );
  NOR2_X1 U443 ( .A1(n580), .A2(n577), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n382), .B(KEYINPUT112), .ZN(n383) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(n383), .ZN(n384) );
  NAND2_X1 U446 ( .A1(n384), .A2(n573), .ZN(n385) );
  NOR2_X1 U447 ( .A1(n555), .A2(n385), .ZN(n386) );
  NOR2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n388), .B(KEYINPUT48), .ZN(n527) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n400) );
  XOR2_X1 U451 ( .A(G211GAT), .B(KEYINPUT21), .Z(n392) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(G218GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n439) );
  XOR2_X1 U454 ( .A(n439), .B(KEYINPUT95), .Z(n394) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(n395), .B(KEYINPUT96), .Z(n398) );
  XNOR2_X1 U458 ( .A(G8GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n515) );
  XNOR2_X1 U461 ( .A(n515), .B(KEYINPUT118), .ZN(n401) );
  NOR2_X1 U462 ( .A1(n527), .A2(n401), .ZN(n402) );
  XNOR2_X1 U463 ( .A(KEYINPUT54), .B(n402), .ZN(n428) );
  XOR2_X1 U464 ( .A(G148GAT), .B(G120GAT), .Z(n404) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(G141GAT), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U467 ( .A(KEYINPUT78), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n427) );
  XOR2_X1 U471 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U474 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n412) );
  XNOR2_X1 U475 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n425) );
  XOR2_X1 U478 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n419), .B(KEYINPUT93), .Z(n423) );
  XOR2_X1 U482 ( .A(G155GAT), .B(KEYINPUT86), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n435), .B(KEYINPUT94), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n513) );
  NAND2_X1 U489 ( .A1(n428), .A2(n513), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n429), .B(KEYINPUT65), .ZN(n567) );
  XOR2_X1 U491 ( .A(G204GAT), .B(KEYINPUT87), .Z(n431) );
  XNOR2_X1 U492 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n446) );
  XOR2_X1 U494 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n433) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U497 ( .A(n434), .B(KEYINPUT85), .Z(n438) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U503 ( .A(n446), .B(n445), .Z(n464) );
  AND2_X1 U504 ( .A1(n567), .A2(n464), .ZN(n449) );
  INV_X1 U505 ( .A(KEYINPUT55), .ZN(n447) );
  NOR2_X1 U506 ( .A1(n519), .A2(n450), .ZN(n563) );
  NAND2_X1 U507 ( .A1(n536), .A2(n563), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n452) );
  XNOR2_X1 U509 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U511 ( .A1(n536), .A2(n577), .ZN(n456) );
  XNOR2_X1 U512 ( .A(KEYINPUT16), .B(n456), .ZN(n473) );
  XOR2_X1 U513 ( .A(n464), .B(KEYINPUT28), .Z(n481) );
  XOR2_X1 U514 ( .A(n515), .B(KEYINPUT27), .Z(n462) );
  INV_X1 U515 ( .A(n462), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n457), .A2(n513), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT97), .ZN(n541) );
  NOR2_X1 U518 ( .A1(n481), .A2(n541), .ZN(n529) );
  XNOR2_X1 U519 ( .A(n529), .B(KEYINPUT98), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n519), .B(KEYINPUT84), .ZN(n459) );
  NAND2_X1 U521 ( .A1(n460), .A2(n459), .ZN(n472) );
  INV_X1 U522 ( .A(n519), .ZN(n528) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(n461), .ZN(n566) );
  NAND2_X1 U524 ( .A1(n566), .A2(n462), .ZN(n467) );
  OR2_X1 U525 ( .A1(n519), .A2(n515), .ZN(n463) );
  NAND2_X1 U526 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n468), .A2(n513), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n473), .A2(n486), .ZN(n474) );
  XOR2_X1 U531 ( .A(n474), .B(KEYINPUT100), .Z(n501) );
  AND2_X1 U532 ( .A1(n573), .A2(n555), .ZN(n490) );
  NAND2_X1 U533 ( .A1(n501), .A2(n490), .ZN(n482) );
  NOR2_X1 U534 ( .A1(n513), .A2(n482), .ZN(n475) );
  XOR2_X1 U535 ( .A(n475), .B(KEYINPUT34), .Z(n476) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  BUF_X1 U537 ( .A(n515), .Z(n504) );
  NOR2_X1 U538 ( .A1(n504), .A2(n482), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(G1325GAT) );
  NOR2_X1 U541 ( .A1(n519), .A2(n482), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n481), .ZN(n523) );
  NOR2_X1 U545 ( .A1(n523), .A2(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n577), .A2(n486), .ZN(n487) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n488) );
  XOR2_X1 U552 ( .A(n489), .B(n488), .Z(n511) );
  AND2_X1 U553 ( .A1(n511), .A2(n490), .ZN(n491) );
  NOR2_X1 U554 ( .A1(n513), .A2(n497), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n497), .A2(n504), .ZN(n494) );
  XOR2_X1 U557 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U558 ( .A1(n519), .A2(n497), .ZN(n495) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(n495), .Z(n496) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n497), .A2(n523), .ZN(n498) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  INV_X1 U563 ( .A(n499), .ZN(n558) );
  NAND2_X1 U564 ( .A1(n558), .A2(n568), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT105), .ZN(n512) );
  NAND2_X1 U566 ( .A1(n512), .A2(n501), .ZN(n507) );
  NOR2_X1 U567 ( .A1(n513), .A2(n507), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(n502), .Z(n503) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n504), .A2(n507), .ZN(n505) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n519), .A2(n507), .ZN(n506) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n523), .A2(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n513), .A2(n522), .ZN(n514) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n522), .ZN(n517) );
  XNOR2_X1 U582 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n522), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U591 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n527), .A2(n530), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n555), .A2(n537), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U597 ( .A1(n537), .A2(n558), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n562), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  NOR2_X1 U606 ( .A1(n527), .A2(n541), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n542), .A2(n566), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n568), .A2(n551), .ZN(n543) );
  XOR2_X1 U609 ( .A(KEYINPUT114), .B(n543), .Z(n544) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  NOR2_X1 U611 ( .A1(n499), .A2(n551), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(KEYINPUT52), .B(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n577), .A2(n551), .ZN(n550) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n563), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  NAND2_X1 U626 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n579), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n579), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

