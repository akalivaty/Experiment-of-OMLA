//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(KEYINPUT74), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(KEYINPUT74), .B2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n208), .A2(new_n210), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n204), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n209), .A2(KEYINPUT75), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G141gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT76), .A4(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n208), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT75), .B(G141gat), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT76), .B1(new_n224), .B2(G148gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n215), .B(new_n218), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n221), .A3(G148gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(new_n222), .A3(new_n208), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n215), .B1(new_n231), .B2(new_n218), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n214), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G113gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT69), .B(G113gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G134gat), .ZN(new_n240));
  INV_X1    g039(.A(G134gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G127gat), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  OAI221_X1 g046(.A(new_n246), .B1(new_n245), .B2(new_n240), .C1(KEYINPUT1), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT70), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n233), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n256), .A2(KEYINPUT82), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(KEYINPUT82), .ZN(new_n258));
  INV_X1    g057(.A(new_n249), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n214), .B(new_n259), .C1(new_n227), .C2(new_n232), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n266), .B(new_n214), .C1(new_n227), .C2(new_n232), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n249), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n263), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n255), .B1(new_n233), .B2(new_n253), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n218), .B1(new_n223), .B2(new_n225), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT77), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n213), .B1(new_n273), .B2(new_n226), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n259), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n270), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n233), .A2(new_n249), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n263), .B1(new_n279), .B2(new_n260), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n280), .B2(new_n264), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n274), .A2(new_n259), .ZN(new_n282));
  AOI211_X1 g081(.A(new_n213), .B(new_n249), .C1(new_n273), .C2(new_n226), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n270), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n264), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT80), .A3(new_n285), .ZN(new_n286));
  AOI221_X4 g085(.A(KEYINPUT81), .B1(new_n277), .B2(new_n268), .C1(new_n281), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n281), .A2(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n277), .A2(new_n268), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n269), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT0), .ZN(new_n294));
  XNOR2_X1  g093(.A(G57gat), .B(G85gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n296), .B(new_n269), .C1(new_n287), .C2(new_n291), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT83), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n292), .A2(new_n297), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT22), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G211gat), .B(G218gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n314), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT27), .B(G183gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n331));
  INV_X1    g130(.A(G183gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(KEYINPUT27), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n329), .ZN(new_n334));
  INV_X1    g133(.A(new_n328), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(KEYINPUT66), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n330), .B1(new_n336), .B2(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G169gat), .ZN(new_n339));
  INV_X1    g138(.A(G176gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT23), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n322), .B2(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT24), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n320), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n342), .B(new_n344), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT64), .B(G176gat), .Z(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT23), .A3(new_n339), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n320), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n346), .B2(new_n320), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n352), .A2(new_n355), .A3(new_n342), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n350), .B1(new_n356), .B2(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G226gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n338), .A2(new_n357), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT29), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n319), .B(new_n362), .C1(new_n364), .C2(new_n361), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n364), .B2(new_n361), .ZN(new_n368));
  OAI221_X1 g167(.A(KEYINPUT73), .B1(new_n359), .B2(new_n360), .C1(new_n363), .C2(KEYINPUT29), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n362), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n370), .B2(new_n318), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT30), .ZN(new_n377));
  INV_X1    g176(.A(new_n371), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n374), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n371), .B2(new_n375), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n202), .B1(new_n308), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT31), .B(G50gat), .Z(new_n384));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n267), .A2(KEYINPUT86), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT86), .B1(new_n267), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n318), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G228gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n266), .B1(new_n318), .B2(KEYINPUT29), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n389), .B(new_n360), .C1(new_n390), .C2(new_n233), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(KEYINPUT87), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n314), .B2(new_n315), .ZN(new_n394));
  INV_X1    g193(.A(new_n314), .ZN(new_n395));
  INV_X1    g194(.A(new_n315), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n314), .A2(new_n393), .A3(new_n315), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n385), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n274), .B1(new_n399), .B2(new_n266), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n319), .B1(new_n267), .B2(new_n385), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n400), .A2(new_n401), .B1(new_n389), .B2(new_n360), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT87), .B1(new_n388), .B2(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(G22gat), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n404), .ZN(new_n406));
  INV_X1    g205(.A(G22gat), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n392), .A4(new_n402), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n405), .B2(new_n408), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n384), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(new_n409), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(new_n384), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n253), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(new_n358), .ZN(new_n420));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n422), .B(KEYINPUT34), .Z(new_n423));
  OR2_X1    g222(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G15gat), .B(G43gat), .Z(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n424), .B(KEYINPUT32), .C1(new_n426), .C2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n423), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n423), .B1(new_n431), .B2(new_n433), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n412), .A2(new_n418), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n304), .B1(new_n300), .B2(new_n301), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n307), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n298), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n379), .A2(new_n381), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(KEYINPUT30), .B2(new_n376), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(KEYINPUT84), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n383), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n307), .A2(new_n301), .A3(new_n300), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n382), .B1(new_n449), .B2(new_n298), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n438), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n289), .A2(new_n290), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n289), .A2(new_n288), .A3(new_n290), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n296), .B1(new_n455), .B2(new_n269), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n298), .B1(new_n302), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n444), .A3(new_n448), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n447), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n444), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n437), .B1(new_n462), .B2(KEYINPUT88), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT35), .B1(new_n450), .B2(new_n448), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT89), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n446), .A2(KEYINPUT35), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n412), .A2(new_n418), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT84), .B1(new_n442), .B2(new_n444), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n202), .B(new_n382), .C1(new_n441), .C2(new_n298), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n436), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n436), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n412), .A2(new_n418), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n262), .A2(new_n268), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n270), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n282), .A2(new_n283), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n263), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n297), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(KEYINPUT39), .B2(new_n479), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n483), .B(KEYINPUT40), .C1(KEYINPUT39), .C2(new_n479), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n307), .A3(new_n382), .A4(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n477), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n378), .A2(KEYINPUT37), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n375), .B1(new_n371), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n370), .A2(new_n319), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n362), .B1(new_n364), .B2(new_n361), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n495), .B(KEYINPUT37), .C1(new_n319), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n376), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n457), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n476), .B1(new_n489), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n470), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n466), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G183gat), .B(G211gat), .Z(new_n504));
  INV_X1    g303(.A(G71gat), .ZN(new_n505));
  INV_X1    g304(.A(G78gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G57gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(G64gat), .ZN(new_n512));
  INV_X1    g311(.A(G64gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(G57gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT9), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n510), .B(new_n515), .C1(new_n508), .C2(new_n509), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(KEYINPUT99), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n512), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n511), .A2(KEYINPUT99), .A3(G64gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n509), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n518), .A2(new_n519), .B1(new_n507), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT100), .Z(new_n523));
  OAI21_X1  g322(.A(new_n516), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT101), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G127gat), .B(G155gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(G1gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT96), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT94), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G1gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n534), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n543), .A2(new_n544), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n537), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G8gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT97), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n525), .B2(new_n524), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n533), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n533), .A2(new_n553), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n504), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  INV_X1    g357(.A(new_n504), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G29gat), .A2(G36gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR3_X1   g364(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G43gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(G50gat), .ZN(new_n569));
  INV_X1    g368(.A(G50gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(G43gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n569), .B2(new_n571), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT15), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(KEYINPUT93), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n568), .B2(G50gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n576), .B(new_n578), .C1(G43gat), .C2(new_n570), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT15), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n567), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n567), .B2(new_n575), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT17), .ZN(new_n584));
  AND3_X1   g383(.A1(KEYINPUT103), .A2(G99gat), .A3(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT103), .B1(G99gat), .B2(G106gat), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT8), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n587), .B(new_n590), .C1(new_n591), .C2(new_n589), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  AND2_X1   g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n596), .A2(new_n583), .B1(KEYINPUT41), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G134gat), .B(G162gat), .Z(new_n604));
  NOR2_X1   g403(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n603), .A2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n562), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n551), .A2(new_n583), .B1(new_n584), .B2(new_n550), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n613), .A2(KEYINPUT18), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(KEYINPUT18), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n551), .B(new_n583), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n612), .B(KEYINPUT13), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G169gat), .B(G197gat), .Z(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT91), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n614), .A2(new_n615), .A3(new_n618), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G230gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n360), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n524), .A2(KEYINPUT104), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n524), .A2(KEYINPUT104), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n634), .A2(new_n635), .A3(new_n594), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n594), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT10), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n594), .A2(new_n639), .A3(new_n524), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT105), .Z(new_n641));
  OAI21_X1  g440(.A(new_n633), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n632), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n503), .A2(new_n610), .A3(new_n630), .A4(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n308), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n382), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n657), .B2(new_n549), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  MUX2_X1   g459(.A(KEYINPUT42), .B(new_n658), .S(new_n660), .Z(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n662), .A3(new_n436), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n653), .A2(new_n476), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n665), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n653), .A2(new_n467), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  OAI21_X1  g468(.A(new_n609), .B1(new_n466), .B2(new_n502), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n630), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n561), .A2(new_n672), .A3(new_n650), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(G29gat), .A3(new_n442), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  OAI211_X1 g475(.A(KEYINPUT106), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n501), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n383), .A2(new_n445), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT106), .B1(new_n679), .B2(new_n467), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n468), .A2(new_n469), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n459), .B1(new_n681), .B2(new_n438), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n448), .B1(new_n457), .B2(new_n444), .ZN(new_n683));
  NOR4_X1   g482(.A1(new_n460), .A2(new_n683), .A3(new_n447), .A4(new_n437), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT89), .B1(new_n463), .B2(new_n464), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI22_X1  g485(.A1(new_n678), .A2(new_n680), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .A4(new_n609), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n670), .A2(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n609), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n470), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n501), .A3(new_n677), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n685), .B2(new_n684), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n693), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n688), .B1(new_n699), .B2(new_n689), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n673), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n442), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n676), .A2(new_n703), .ZN(G1328gat));
  INV_X1    g503(.A(G36gat), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n671), .A2(new_n705), .A3(new_n382), .A4(new_n673), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  OAI211_X1 g506(.A(new_n382), .B(new_n673), .C1(new_n692), .C2(new_n700), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G36gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(KEYINPUT108), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(new_n436), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n568), .B1(new_n674), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n476), .A2(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n702), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n720), .B(new_n716), .C1(new_n702), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1330gat));
  NOR3_X1   g521(.A1(new_n674), .A2(G50gat), .A3(new_n477), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n467), .B(new_n673), .C1(new_n692), .C2(new_n700), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(G50gat), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT109), .B1(new_n724), .B2(G50gat), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI221_X4 g527(.A(new_n723), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n724), .C2(G50gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  AND4_X1   g529(.A1(new_n610), .A2(new_n687), .A3(new_n672), .A4(new_n650), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n308), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n382), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT110), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT111), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n735), .B(new_n738), .ZN(G1333gat));
  AOI21_X1  g538(.A(new_n505), .B1(new_n731), .B2(new_n476), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n436), .B(KEYINPUT112), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G71gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n731), .A2(new_n467), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g546(.A1(new_n561), .A2(new_n630), .A3(new_n651), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n308), .B(new_n748), .C1(new_n692), .C2(new_n700), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G85gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n442), .A2(G85gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n561), .A2(new_n630), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n699), .B2(new_n752), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n650), .B(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1336gat));
  OAI211_X1 g557(.A(new_n382), .B(new_n748), .C1(new_n692), .C2(new_n700), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n444), .A2(G92gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n650), .B(new_n762), .C1(new_n753), .C2(new_n754), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g564(.A1(new_n701), .A2(new_n476), .A3(new_n748), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G99gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n715), .A2(new_n651), .A3(G99gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n753), .B2(new_n754), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1338gat));
  OAI211_X1 g569(.A(new_n467), .B(new_n748), .C1(new_n692), .C2(new_n700), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n477), .A2(G106gat), .A3(new_n651), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n753), .B2(new_n754), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n774), .B2(KEYINPUT115), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n775), .B(new_n777), .ZN(G1339gat));
  OR3_X1    g577(.A1(new_n638), .A2(new_n641), .A3(new_n633), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(KEYINPUT54), .A3(new_n642), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(new_n633), .C1(new_n638), .C2(new_n641), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n782), .A2(new_n783), .A3(new_n647), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n782), .B2(new_n647), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(KEYINPUT55), .B(new_n780), .C1(new_n784), .C2(new_n785), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n630), .A2(new_n648), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT117), .B1(new_n611), .B2(new_n612), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n616), .B2(new_n617), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n611), .A2(KEYINPUT117), .A3(new_n612), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n625), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n629), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n650), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n609), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n609), .ZN(new_n799));
  INV_X1    g598(.A(new_n788), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n789), .A2(new_n648), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n803), .A3(KEYINPUT118), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n797), .B2(new_n802), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n561), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n561), .A2(new_n693), .A3(new_n672), .A4(new_n651), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(new_n442), .A3(new_n382), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n438), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n811), .A2(new_n236), .A3(new_n672), .ZN(new_n812));
  INV_X1    g611(.A(new_n809), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT119), .A3(new_n477), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n809), .B2(new_n467), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n442), .A2(new_n382), .A3(new_n715), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n817), .A2(KEYINPUT120), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT120), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n672), .ZN(new_n821));
  INV_X1    g620(.A(G113gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n812), .B1(new_n821), .B2(new_n822), .ZN(G1340gat));
  INV_X1    g622(.A(new_n811), .ZN(new_n824));
  AOI21_X1  g623(.A(G120gat), .B1(new_n824), .B2(new_n650), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n819), .A2(new_n820), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n651), .A2(new_n234), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(G1341gat));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n239), .A3(new_n561), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n819), .A2(new_n820), .A3(new_n562), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n239), .ZN(G1342gat));
  NAND4_X1  g630(.A1(new_n810), .A2(new_n241), .A3(new_n438), .A4(new_n609), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT56), .Z(new_n833));
  NOR3_X1   g632(.A1(new_n819), .A2(new_n820), .A3(new_n693), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n241), .ZN(G1343gat));
  NOR2_X1   g634(.A1(new_n442), .A2(new_n382), .ZN(new_n836));
  INV_X1    g635(.A(new_n476), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n561), .B1(new_n798), .B2(new_n803), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n467), .B1(new_n839), .B2(new_n808), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n842), .B(new_n467), .C1(new_n807), .C2(new_n808), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n843), .A3(new_n630), .ZN(new_n844));
  INV_X1    g643(.A(new_n224), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n476), .A2(new_n477), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n836), .B(new_n846), .C1(new_n807), .C2(new_n808), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n672), .A2(G141gat), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n844), .A2(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT122), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n850), .B2(new_n851), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n853), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n853), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n207), .A2(KEYINPUT59), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n848), .B2(new_n650), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n813), .A2(KEYINPUT57), .A3(new_n467), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n840), .A2(new_n842), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n650), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n836), .A2(KEYINPUT59), .A3(new_n837), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n843), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n651), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n866), .A2(new_n867), .B1(KEYINPUT59), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n862), .B1(new_n870), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g670(.A(G155gat), .B1(new_n868), .B2(new_n562), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n562), .A2(G155gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n847), .B2(new_n873), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n868), .B2(new_n693), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n693), .A2(G162gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n847), .B2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n809), .A2(new_n308), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n437), .A2(new_n444), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(G169gat), .B1(new_n881), .B2(new_n630), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n442), .A2(new_n382), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT123), .Z(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n741), .B(new_n885), .C1(new_n814), .C2(new_n816), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n672), .A2(new_n339), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n881), .B2(new_n650), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n651), .A2(new_n351), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n886), .B2(new_n890), .ZN(G1349gat));
  NAND2_X1  g690(.A1(new_n561), .A2(new_n328), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n881), .A2(KEYINPUT124), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n880), .B2(new_n892), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n885), .A2(new_n741), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n817), .A2(new_n561), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n897), .B(new_n898), .C1(new_n332), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n332), .B1(new_n886), .B2(new_n561), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n894), .A2(new_n896), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT60), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n881), .A2(new_n329), .A3(new_n609), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n886), .A2(new_n609), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(G190gat), .ZN(new_n909));
  AOI211_X1 g708(.A(KEYINPUT61), .B(new_n329), .C1(new_n886), .C2(new_n609), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(G1351gat));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n885), .A2(new_n476), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n865), .A2(new_n630), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(KEYINPUT125), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(KEYINPUT125), .B2(new_n914), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n476), .A2(new_n444), .A3(new_n477), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n878), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n912), .A3(new_n630), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(G1352gat));
  NOR3_X1   g720(.A1(new_n918), .A2(G204gat), .A3(new_n651), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  INV_X1    g722(.A(G204gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n866), .A2(new_n476), .A3(new_n885), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n309), .A3(new_n561), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n865), .A2(new_n561), .A3(new_n913), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(new_n310), .B1(new_n918), .B2(new_n693), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n865), .A2(G218gat), .A3(new_n609), .A4(new_n913), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT126), .B(new_n310), .C1(new_n918), .C2(new_n693), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


