//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  XOR2_X1   g000(.A(KEYINPUT71), .B(G902), .Z(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G140), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT16), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n189), .B2(KEYINPUT16), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT74), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n199), .A3(G146), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n189), .A2(new_n191), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n209), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n198), .A2(new_n200), .A3(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n192), .C1(new_n193), .C2(new_n195), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n197), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(new_n208), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n211), .A2(new_n212), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT65), .A2(G953), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT65), .A2(G953), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n229));
  AND2_X1   g043(.A1(G221), .A2(G234), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n228), .B2(new_n230), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n225), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n233), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n231), .A3(new_n224), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n217), .A2(new_n223), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n217), .A2(new_n223), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT76), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT76), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n187), .B(new_n238), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n217), .A2(new_n223), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n242), .A3(new_n241), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n246), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n249), .A2(new_n187), .A3(new_n238), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G217), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n187), .B2(G234), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G902), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n249), .A2(new_n238), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n252), .A2(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  NOR2_X1   g073(.A1(G472), .A2(G902), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n228), .A2(G210), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT26), .B(G101), .Z(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n268), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT2), .B(G113), .Z(new_n274));
  OR2_X1    g088(.A1(KEYINPUT64), .A2(G116), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT64), .A2(G116), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(G119), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n202), .A2(G116), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n278), .B2(new_n277), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  INV_X1    g099(.A(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT11), .A3(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(G137), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G131), .ZN(new_n290));
  INV_X1    g104(.A(G131), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n285), .A2(new_n287), .A3(new_n291), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n214), .A2(G143), .ZN(new_n294));
  INV_X1    g108(.A(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G146), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G143), .B(G146), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT0), .B(G128), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT1), .B1(new_n295), .B2(G146), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n295), .A2(G146), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n214), .A2(G143), .ZN(new_n306));
  OAI211_X1 g120(.A(G128), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n284), .A2(G137), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n286), .A2(G134), .ZN(new_n309));
  OAI21_X1  g123(.A(G131), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n294), .B(new_n296), .C1(KEYINPUT1), .C2(new_n205), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n307), .A2(new_n292), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n282), .A2(new_n303), .A3(KEYINPUT28), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n281), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n279), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n301), .B1(new_n292), .B2(new_n290), .ZN(new_n316));
  INV_X1    g130(.A(new_n312), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n282), .A2(new_n303), .A3(new_n312), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n273), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT30), .B1(new_n316), .B2(new_n317), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n303), .A2(new_n327), .A3(new_n312), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n329), .B2(new_n315), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT31), .B1(new_n330), .B2(new_n273), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n282), .B1(new_n326), .B2(new_n328), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT31), .ZN(new_n333));
  NOR4_X1   g147(.A1(new_n332), .A2(new_n272), .A3(new_n333), .A4(new_n325), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n324), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT67), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT30), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n327), .B1(new_n303), .B2(new_n312), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n315), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n273), .A3(new_n320), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n333), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n273), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT67), .A3(new_n324), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n261), .B1(new_n337), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n259), .B1(new_n346), .B2(KEYINPUT32), .ZN(new_n347));
  INV_X1    g161(.A(G472), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT70), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT70), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n315), .B(new_n350), .C1(new_n316), .C2(new_n317), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(KEYINPUT28), .A3(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(KEYINPUT29), .A3(new_n273), .A4(new_n322), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(new_n187), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n319), .A2(new_n273), .A3(new_n322), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT69), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n272), .B1(new_n332), .B2(new_n325), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT69), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n319), .A2(new_n273), .A3(new_n359), .A4(new_n322), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n348), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n346), .B2(KEYINPUT32), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT67), .B1(new_n344), .B2(new_n324), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n336), .B(new_n323), .C1(new_n342), .C2(new_n343), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n260), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT68), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n347), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n363), .A2(new_n347), .A3(new_n368), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n258), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G214), .B1(G237), .B2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G210), .B1(G237), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n315), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n390), .B2(G101), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT78), .B(G107), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n396), .A2(new_n381), .B1(KEYINPUT3), .B2(new_n387), .ZN(new_n397));
  AOI21_X1  g211(.A(G101), .B1(new_n380), .B2(G107), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT79), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n386), .A2(KEYINPUT79), .A3(new_n388), .A4(new_n398), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n386), .A2(new_n388), .A3(new_n398), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n400), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT80), .A3(new_n395), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n394), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n387), .B1(new_n396), .B2(G104), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G101), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n277), .A2(KEYINPUT5), .A3(new_n278), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n202), .A3(G116), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(G113), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n279), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n379), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n282), .B1(new_n392), .B2(new_n391), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n408), .A2(KEYINPUT80), .A3(new_n395), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT80), .B1(new_n408), .B2(new_n395), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n419), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n378), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n301), .A2(G125), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n307), .A2(new_n311), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n430), .B2(G125), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(G224), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G953), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n431), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n379), .C1(new_n410), .C2(new_n419), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(new_n432), .B2(G953), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n431), .B(new_n438), .Z(new_n439));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n378), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n408), .A2(KEYINPUT83), .A3(new_n412), .ZN(new_n443));
  INV_X1    g257(.A(new_n418), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n407), .A2(new_n400), .B1(G101), .B2(new_n411), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n418), .B1(new_n446), .B2(KEYINPUT83), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n440), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(new_n444), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n418), .A3(KEYINPUT83), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n450), .A4(new_n442), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n426), .A2(new_n439), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G902), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n437), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT85), .B1(new_n452), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n377), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n453), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(new_n376), .A3(new_n437), .A4(new_n454), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n375), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G221), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT9), .B(G234), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n463), .B1(new_n465), .B2(new_n453), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n228), .A2(G227), .ZN(new_n467));
  XOR2_X1   g281(.A(G110), .B(G140), .Z(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n446), .A2(new_n430), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n408), .A2(new_n430), .A3(new_n412), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n293), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n293), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n413), .A2(new_n429), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n408), .A2(new_n430), .A3(new_n412), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT12), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n301), .B1(new_n391), .B2(new_n392), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n422), .B2(new_n423), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(KEYINPUT10), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT10), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n446), .A2(new_n485), .A3(new_n430), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n487), .A3(new_n476), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n470), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n483), .A2(new_n487), .A3(new_n476), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n476), .B1(new_n483), .B2(new_n487), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n490), .A2(new_n491), .A3(new_n469), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G469), .B1(new_n493), .B2(G902), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n469), .B1(new_n490), .B2(new_n491), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n479), .A2(KEYINPUT12), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n488), .B(new_n470), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n187), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n466), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n295), .A2(G128), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(KEYINPUT91), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n205), .B2(G143), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n295), .A2(KEYINPUT90), .A3(G128), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n504), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n506), .A2(new_n510), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G134), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n284), .B(new_n504), .C1(new_n508), .C2(new_n509), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n275), .A2(G122), .A3(new_n276), .ZN(new_n518));
  INV_X1    g332(.A(G122), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G116), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n396), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n396), .A3(new_n520), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(KEYINPUT88), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n525));
  INV_X1    g339(.A(new_n523), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(new_n521), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n516), .A2(new_n517), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G134), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n530), .B2(new_n517), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n520), .B1(new_n518), .B2(KEYINPUT14), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n518), .A2(KEYINPUT14), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n518), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n537), .B2(new_n382), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n464), .A2(new_n253), .A3(G953), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n528), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n528), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n187), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT93), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n187), .C1(new_n540), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n542), .B2(KEYINPUT93), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n553));
  INV_X1    g367(.A(new_n227), .ZN(new_n554));
  NAND2_X1  g368(.A1(KEYINPUT65), .A2(G953), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n554), .A2(G214), .A3(new_n262), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n295), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n228), .A2(G143), .A3(G214), .A4(new_n262), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n553), .B(new_n291), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT87), .B1(new_n219), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT17), .A3(G131), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n218), .A4(new_n197), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(G131), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n557), .A2(new_n558), .A3(new_n291), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n553), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n561), .A2(KEYINPUT18), .A3(G131), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n215), .B(new_n214), .ZN(new_n570));
  NAND2_X1  g384(.A1(KEYINPUT18), .A2(G131), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n557), .A2(new_n558), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G113), .B(G122), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT86), .B(G104), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n568), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n568), .B2(new_n573), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n453), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G475), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT20), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n568), .A2(new_n573), .A3(new_n577), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n565), .A2(new_n566), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n215), .B(KEYINPUT19), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n214), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n584), .A2(new_n198), .A3(new_n200), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n573), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n576), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G475), .A2(G902), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT20), .B(new_n593), .C1(new_n583), .C2(new_n589), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n581), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G953), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G952), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(G234), .B2(G237), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT21), .B(G898), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT94), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n228), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n552), .A2(new_n595), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n462), .A2(new_n502), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n373), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(new_n466), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n483), .A2(new_n487), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n293), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n488), .A3(new_n470), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n483), .A2(new_n487), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n476), .A2(new_n612), .B1(new_n475), .B2(new_n480), .ZN(new_n613));
  OAI211_X1 g427(.A(G469), .B(new_n611), .C1(new_n613), .C2(new_n470), .ZN(new_n614));
  NAND2_X1  g428(.A1(G469), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n187), .ZN(new_n617));
  AOI211_X1 g431(.A(G469), .B(new_n617), .C1(new_n495), .C2(new_n498), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n257), .B(new_n608), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n337), .B2(new_n345), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n366), .B1(new_n620), .B2(new_n348), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n542), .A2(new_n547), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n540), .A2(new_n541), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT95), .B1(new_n528), .B2(new_n538), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n187), .A2(G478), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n595), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n457), .A2(new_n461), .ZN(new_n635));
  INV_X1    g449(.A(new_n603), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n374), .A3(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n623), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND2_X1  g454(.A1(new_n590), .A2(new_n591), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT20), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n590), .A2(new_n582), .A3(new_n591), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(KEYINPUT96), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n592), .B2(new_n594), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n580), .A2(new_n648), .A3(G475), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n580), .B2(G475), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(new_n651), .A3(new_n552), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n623), .A2(new_n637), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n252), .A2(new_n254), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT36), .B1(new_n241), .B2(new_n242), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n248), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n255), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n660), .B(new_n608), .C1(new_n616), .C2(new_n618), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n621), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n462), .A3(new_n604), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  NAND3_X1  g479(.A1(new_n462), .A2(new_n502), .A3(new_n660), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n370), .B2(new_n372), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n598), .B1(new_n602), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n652), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(new_n669), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n502), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n502), .A2(KEYINPUT40), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n330), .A2(new_n272), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(G902), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n349), .A2(new_n351), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n272), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n348), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n346), .B2(KEYINPUT32), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n347), .A2(new_n685), .A3(new_n368), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n635), .B(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n552), .A2(new_n595), .A3(new_n374), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n660), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n679), .A2(new_n689), .A3(new_n690), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND2_X1  g510(.A1(new_n370), .A2(new_n372), .ZN(new_n697));
  INV_X1    g511(.A(new_n666), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n634), .B2(new_n669), .ZN(new_n700));
  INV_X1    g514(.A(new_n669), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n633), .A2(new_n595), .A3(KEYINPUT100), .A4(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n697), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  NAND2_X1  g519(.A1(new_n499), .A2(new_n187), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n608), .A3(new_n501), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n637), .A2(new_n634), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n373), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT41), .B(G113), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT101), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n710), .B(new_n712), .ZN(G15));
  NOR3_X1   g527(.A1(new_n637), .A2(new_n652), .A3(new_n708), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n373), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  INV_X1    g530(.A(new_n708), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(new_n462), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n604), .A2(new_n660), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n697), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  AOI21_X1  g535(.A(new_n693), .B1(new_n457), .B2(new_n461), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n352), .A2(new_n322), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n344), .B1(new_n723), .B2(new_n273), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n260), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n257), .B(new_n725), .C1(new_n620), .C2(new_n348), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n722), .A2(new_n636), .A3(new_n717), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT102), .B(G122), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G24));
  NAND2_X1  g544(.A1(new_n700), .A2(new_n702), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n660), .B(new_n725), .C1(new_n620), .C2(new_n348), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n718), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  NAND3_X1  g549(.A1(new_n457), .A2(new_n374), .A3(new_n461), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT103), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n457), .A2(new_n738), .A3(new_n374), .A4(new_n461), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n502), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(KEYINPUT104), .A3(new_n502), .A4(new_n739), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n373), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n366), .A2(new_n367), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n258), .B1(new_n363), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n703), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n742), .B2(new_n743), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n746), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n291), .ZN(G33));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n373), .A3(new_n670), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  AND2_X1   g569(.A1(new_n633), .A2(KEYINPUT43), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n595), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n581), .B(KEYINPUT105), .C1(new_n592), .C2(new_n594), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n756), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n595), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n766), .B2(new_n633), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT44), .A3(new_n621), .A4(new_n660), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n737), .A2(new_n739), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n767), .B1(new_n761), .B2(new_n764), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n621), .A2(new_n660), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n493), .A2(KEYINPUT45), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n489), .B2(new_n492), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(G469), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n615), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n618), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n615), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n466), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(new_n673), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n770), .A2(new_n772), .A3(new_n776), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  OR2_X1    g602(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n793));
  NAND2_X1  g607(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n789), .A2(new_n792), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n797), .B(new_n466), .C1(new_n783), .C2(new_n784), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n790), .B(new_n791), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n697), .A2(new_n257), .A3(new_n731), .A4(new_n771), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  AND2_X1   g617(.A1(new_n707), .A2(new_n501), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT109), .Z(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n608), .A2(new_n762), .A3(new_n374), .A4(new_n633), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n692), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n810), .A2(new_n258), .A3(new_n689), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n744), .A2(new_n733), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n669), .B(new_n550), .C1(new_n546), .C2(new_n548), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n647), .A2(new_n651), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(new_n661), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n771), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n818), .A2(new_n697), .A3(KEYINPUT110), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT110), .B1(new_n818), .B2(new_n697), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n697), .B(new_n257), .C1(new_n709), .C2(new_n714), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n375), .B(new_n603), .C1(new_n457), .C2(new_n461), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n766), .A2(new_n552), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n634), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n622), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n728), .A2(new_n826), .A3(new_n663), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n822), .A2(new_n606), .A3(new_n827), .A4(new_n720), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n744), .A2(new_n373), .A3(new_n670), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n752), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n660), .A2(new_n669), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n722), .A2(new_n686), .A3(new_n502), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n671), .A2(new_n704), .A3(new_n734), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n667), .A2(new_n670), .B1(new_n718), .B2(new_n733), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .A3(new_n704), .A4(new_n833), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n813), .A2(new_n830), .A3(new_n831), .A4(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n754), .B(new_n814), .C1(new_n820), .C2(new_n819), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n752), .A3(new_n828), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n813), .B1(new_n842), .B2(new_n839), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n812), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n830), .A2(new_n831), .A3(new_n839), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n813), .A3(new_n839), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(KEYINPUT112), .A3(new_n812), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n839), .B2(KEYINPUT111), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n847), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n842), .B(new_n839), .C1(KEYINPUT111), .C2(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n805), .A2(new_n466), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n795), .A2(new_n799), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n727), .A2(new_n598), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n774), .A2(new_n771), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n598), .A2(new_n737), .A3(new_n717), .A4(new_n739), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n769), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n732), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n257), .A3(new_n687), .A4(new_n688), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n633), .A2(new_n595), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT116), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  OAI221_X1 g683(.A(new_n869), .B1(new_n865), .B2(new_n866), .C1(new_n732), .C2(new_n863), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n692), .A2(new_n375), .A3(new_n717), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n692), .A2(KEYINPUT114), .A3(new_n375), .A4(new_n717), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n877));
  NOR2_X1   g691(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n774), .A2(new_n859), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n876), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n861), .A2(new_n871), .A3(new_n882), .A4(KEYINPUT51), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n769), .A2(new_n749), .A3(new_n862), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT48), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT118), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n769), .A2(new_n598), .A3(new_n718), .A4(new_n727), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n597), .B(KEYINPUT117), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n888), .B(new_n889), .C1(new_n865), .C2(new_n634), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n887), .B(new_n890), .C1(new_n884), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NOR4_X1   g707(.A1(new_n880), .A2(new_n881), .A3(new_n864), .A4(new_n867), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n857), .B(KEYINPUT113), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n860), .B1(new_n800), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT51), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n846), .A2(new_n851), .A3(new_n856), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT120), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n899), .B2(new_n900), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n811), .B1(new_n901), .B2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n840), .A2(new_n843), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n617), .A3(new_n377), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n427), .A2(new_n436), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n434), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT55), .Z(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n228), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n907), .B2(KEYINPUT121), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(KEYINPUT121), .B2(new_n907), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n917), .B2(new_n910), .ZN(G51));
  XNOR2_X1  g732(.A(new_n850), .B(KEYINPUT54), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n615), .B(KEYINPUT57), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n499), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n850), .A2(new_n187), .A3(new_n780), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(G54));
  NAND4_X1  g737(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .A4(new_n617), .ZN(new_n924));
  INV_X1    g738(.A(new_n590), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n913), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n629), .A2(new_n630), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n914), .B1(new_n919), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n846), .A2(new_n851), .A3(new_n856), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n631), .B2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT122), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n906), .A2(new_n658), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n906), .A2(new_n939), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n914), .B(new_n940), .C1(new_n941), .C2(new_n256), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n601), .B2(new_n432), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT123), .Z(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n828), .B2(new_n228), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n908), .B1(G898), .B2(new_n228), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n947), .B(new_n948), .Z(G69));
  INV_X1    g763(.A(new_n674), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n373), .A2(new_n772), .A3(new_n950), .A4(new_n825), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n787), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n671), .A2(new_n704), .A3(new_n734), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n695), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n695), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n802), .A2(new_n952), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n228), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n329), .B(new_n585), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n228), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n787), .A2(new_n953), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n786), .A2(new_n722), .A3(new_n749), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n752), .A2(new_n966), .A3(new_n829), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n802), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n963), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n228), .A2(G900), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n961), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT124), .ZN(new_n973));
  INV_X1    g787(.A(G227), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n962), .B1(new_n974), .B2(new_n668), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n961), .A2(new_n969), .A3(new_n976), .A4(new_n971), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n975), .B1(new_n973), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  OR2_X1    g796(.A1(new_n965), .A2(new_n968), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n828), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n272), .A3(new_n330), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n958), .B2(new_n828), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n913), .B1(new_n986), .B2(new_n680), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n357), .B(KEYINPUT126), .Z(new_n989));
  INV_X1    g803(.A(new_n341), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n982), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT127), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n855), .B2(new_n992), .ZN(G57));
endmodule


