//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(new_n454), .B2(G2106), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n456), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n454), .A2(KEYINPUT65), .A3(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n465), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n466), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n465), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n475), .A2(G137), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(new_n475), .A2(new_n477), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(KEYINPUT67), .A3(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n476), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n484), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n476), .A3(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n469), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n475), .A2(G138), .A3(new_n476), .A4(new_n477), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  XOR2_X1   g076(.A(KEYINPUT68), .B(G114), .Z(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(new_n476), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n475), .A2(G126), .A3(G2105), .A4(new_n477), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n499), .A2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT69), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT70), .B(G88), .Z(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n508), .A2(G543), .A3(new_n515), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n507), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n521), .A2(G51), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI211_X1 g108(.A(new_n531), .B(new_n532), .C1(new_n513), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n508), .A2(G52), .A3(G543), .A4(new_n515), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n508), .A2(G90), .A3(new_n513), .A4(new_n515), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n541), .A2(KEYINPUT71), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(KEYINPUT71), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n510), .A2(new_n512), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n507), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT72), .ZN(new_n552));
  AOI22_X1  g127(.A1(G43), .A2(new_n521), .B1(new_n517), .B2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT73), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n515), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n547), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n517), .A2(G91), .B1(G651), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n521), .A2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n517), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n513), .A2(G61), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(new_n575), .B1(G73), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n576), .B1(new_n575), .B2(new_n574), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(new_n550), .B1(G48), .B2(new_n521), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n517), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT75), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n517), .A2(new_n581), .A3(G86), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G60), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n547), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(new_n550), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(G47), .A2(new_n521), .B1(new_n517), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n517), .A2(new_n592), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT77), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n547), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n514), .B1(new_n599), .B2(KEYINPUT79), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(KEYINPUT79), .B2(new_n599), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n520), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(new_n520), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n596), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT10), .B1(new_n593), .B2(new_n595), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT80), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  MUX2_X1   g185(.A(G301), .B(new_n609), .S(new_n610), .Z(G284));
  XNOR2_X1  g186(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(new_n609), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT82), .B(G559), .Z(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(G860), .B2(new_n618), .ZN(G148));
  NAND2_X1  g194(.A1(new_n554), .A2(new_n610), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n622), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g199(.A1(new_n483), .A2(KEYINPUT83), .A3(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n486), .A2(G135), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n482), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n625), .A2(new_n626), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(KEYINPUT17), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n657), .A2(new_n655), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n661), .B2(new_n657), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT85), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT86), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(KEYINPUT86), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT21), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G25), .A2(G29), .ZN(new_n695));
  OR2_X1    g270(.A1(G95), .A2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n697));
  INV_X1    g272(.A(G131), .ZN(new_n698));
  INV_X1    g273(.A(G119), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n697), .B1(new_n485), .B2(new_n698), .C1(new_n699), .C2(new_n482), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n695), .B1(new_n701), .B2(G29), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1986), .Z(new_n710));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n711));
  INV_X1    g286(.A(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(G16), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G303), .B2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1971), .ZN(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G23), .ZN(new_n718));
  INV_X1    g293(.A(G288), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT33), .B(G1976), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  AND2_X1   g297(.A1(new_n706), .A2(G6), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G305), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n717), .A2(new_n722), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n705), .B(new_n710), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n617), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1348), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n706), .A2(G20), .ZN(new_n737));
  OAI211_X1 g312(.A(KEYINPUT23), .B(new_n737), .C1(new_n614), .C2(new_n706), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT23), .B2(new_n737), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n742), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT94), .Z(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G35), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G162), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2090), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n740), .B1(new_n741), .B2(new_n746), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n742), .A2(G26), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n483), .A2(G128), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n486), .A2(G140), .ZN(new_n756));
  OR2_X1    g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n742), .ZN(new_n761));
  MUX2_X1   g336(.A(new_n754), .B(new_n761), .S(KEYINPUT28), .Z(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G2067), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n706), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n706), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(G2067), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n742), .A2(G33), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n472), .A2(G103), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n486), .B2(G139), .ZN(new_n773));
  NAND2_X1  g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  INV_X1    g349(.A(G127), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n469), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n476), .B1(new_n777), .B2(KEYINPUT93), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(KEYINPUT93), .B2(new_n777), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n769), .B1(new_n780), .B2(new_n742), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2072), .ZN(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G32), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT26), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(G105), .B2(new_n472), .ZN(new_n788));
  INV_X1    g363(.A(G141), .ZN(new_n789));
  INV_X1    g364(.A(G129), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n788), .B1(new_n485), .B2(new_n789), .C1(new_n790), .C2(new_n482), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n783), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT27), .B(G1996), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n706), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n706), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1966), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n782), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n742), .B1(KEYINPUT24), .B2(G34), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(KEYINPUT24), .B2(G34), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n479), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2084), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT30), .B(G28), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n804), .A2(new_n742), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n803), .B(new_n807), .C1(new_n742), .C2(new_n632), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n706), .A2(G19), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n555), .B2(new_n706), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1341), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n808), .B(new_n811), .C1(G1961), .C2(new_n765), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n751), .A2(new_n752), .B1(new_n741), .B2(new_n746), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n768), .A2(new_n799), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n733), .A2(new_n736), .A3(new_n753), .A4(new_n814), .ZN(G311));
  OR4_X1    g390(.A1(new_n733), .A2(new_n736), .A3(new_n753), .A4(new_n814), .ZN(G150));
  NAND2_X1  g391(.A1(new_n517), .A2(G93), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n521), .A2(G55), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n507), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  INV_X1    g397(.A(G559), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT39), .B1(new_n609), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n609), .A2(KEYINPUT39), .A3(new_n823), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT96), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n826), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(new_n829), .A3(new_n824), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n554), .B(new_n820), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n827), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n833), .ZN(new_n839));
  INV_X1    g414(.A(new_n835), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n834), .B1(new_n827), .B2(new_n830), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT97), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  AND4_X1   g418(.A1(KEYINPUT97), .A2(new_n842), .A3(new_n836), .A4(new_n837), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n822), .B1(new_n843), .B2(new_n844), .ZN(G145));
  XOR2_X1   g420(.A(new_n700), .B(new_n791), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n780), .ZN(new_n847));
  INV_X1    g422(.A(new_n505), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n849));
  INV_X1    g424(.A(new_n497), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT99), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n852));
  AOI211_X1 g427(.A(new_n852), .B(new_n497), .C1(new_n498), .C2(KEYINPUT4), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n759), .B(new_n854), .Z(new_n855));
  OR2_X1    g430(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n847), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n483), .A2(G130), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n486), .A2(G142), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n476), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n635), .B(KEYINPUT100), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n479), .B(KEYINPUT98), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n493), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n632), .Z(new_n870));
  NAND3_X1  g445(.A1(new_n856), .A2(new_n865), .A3(new_n857), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT101), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n867), .A2(new_n875), .A3(new_n870), .A4(new_n871), .ZN(new_n876));
  INV_X1    g451(.A(new_n870), .ZN(new_n877));
  INV_X1    g452(.A(new_n871), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n865), .B1(new_n856), .B2(new_n857), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n873), .A2(new_n874), .A3(new_n876), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(G395));
  NAND2_X1  g458(.A1(new_n622), .A2(new_n833), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n621), .A2(new_n839), .ZN(new_n885));
  NAND2_X1  g460(.A1(G299), .A2(KEYINPUT103), .ZN(new_n886));
  OR2_X1    g461(.A1(G299), .A2(KEYINPUT103), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n608), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(KEYINPUT103), .B(G299), .C1(new_n606), .C2(new_n607), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n621), .B(new_n833), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT41), .B1(new_n888), .B2(new_n889), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n891), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND2_X1  g473(.A1(G305), .A2(G290), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n580), .A2(new_n582), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n708), .A2(new_n900), .A3(new_n578), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(G288), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G288), .B1(new_n899), .B2(new_n901), .ZN(new_n904));
  XOR2_X1   g479(.A(G303), .B(KEYINPUT104), .Z(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n719), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n909), .B2(new_n902), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n898), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n906), .B1(new_n903), .B2(new_n904), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n905), .A3(new_n902), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n907), .B2(new_n910), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n897), .A2(new_n916), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n916), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n897), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n897), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n820), .A2(new_n610), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(new_n538), .C1(new_n542), .C2(new_n543), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(G168), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G168), .B1(new_n930), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n839), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G286), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n833), .A3(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n895), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n939), .A3(KEYINPUT108), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n943), .B(new_n839), .C1(new_n934), .C2(new_n935), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n890), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n915), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n947), .A2(new_n874), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n941), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n907), .A2(new_n910), .A3(new_n898), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT105), .B1(new_n912), .B2(new_n913), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n929), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n936), .A2(new_n939), .A3(new_n890), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n945), .B2(new_n896), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n947), .A3(new_n874), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n928), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n928), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n948), .A2(new_n929), .A3(new_n953), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT109), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT109), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G397));
  XOR2_X1   g540(.A(KEYINPUT110), .B(G1384), .Z(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n854), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n471), .A2(G2105), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n472), .A2(G101), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(G40), .A3(new_n478), .A4(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n473), .A2(KEYINPUT111), .A3(G40), .A4(new_n478), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n791), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(G1996), .B2(new_n975), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(G1996), .B2(new_n792), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n759), .B(G2067), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT113), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n700), .B(new_n703), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n975), .ZN(new_n987));
  XNOR2_X1  g562(.A(G290), .B(G1986), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n854), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n499), .B2(new_n505), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n972), .A2(new_n973), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n990), .B1(new_n996), .B2(G2078), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n854), .A2(new_n992), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n994), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n974), .C1(new_n994), .C2(new_n993), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n741), .A2(KEYINPUT53), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n993), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT115), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n974), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n854), .A2(new_n1005), .A3(new_n992), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n854), .A2(new_n1008), .A3(new_n1005), .A4(new_n992), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1004), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g585(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .C1(new_n1010), .C2(G1961), .ZN(new_n1011));
  XNOR2_X1  g586(.A(G301), .B(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n967), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n970), .A2(new_n1001), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n991), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1012), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(new_n997), .C1(G1961), .C2(new_n1010), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  INV_X1    g595(.A(G2084), .ZN(new_n1021));
  INV_X1    g596(.A(G1966), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1010), .A2(new_n1021), .B1(new_n1000), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(G168), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G168), .A2(new_n1020), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1000), .A2(new_n1022), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1024), .A2(new_n1025), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1026), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT51), .B(new_n1031), .C1(new_n1023), .C2(new_n1020), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1019), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n974), .A2(new_n854), .A3(new_n992), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n578), .A2(new_n579), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G1981), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n900), .A2(new_n1038), .A3(new_n578), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1035), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1034), .B(G8), .C1(new_n1044), .C2(G288), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n719), .A2(G1976), .ZN(new_n1046));
  OR3_X1    g621(.A1(new_n1045), .A2(KEYINPUT52), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1971), .B1(new_n991), .B2(new_n995), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1004), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n752), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1053), .B2(KEYINPUT116), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1010), .A2(new_n1055), .A3(new_n752), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1020), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND4_X1  g637(.A1(G303), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT118), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1049), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1005), .B1(new_n854), .B2(new_n992), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n974), .B1(KEYINPUT50), .B2(new_n993), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1067), .A2(new_n1068), .A3(G2090), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1069), .B2(new_n1050), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1064), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT125), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1053), .A2(KEYINPUT116), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1050), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n1056), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(G8), .A3(new_n1065), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1049), .ZN(new_n1077));
  AND4_X1   g652(.A1(KEYINPUT125), .A2(new_n1076), .A3(new_n1071), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1033), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1956), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n991), .A2(new_n995), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(G299), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  AOI211_X1 g662(.A(KEYINPUT120), .B(new_n1087), .C1(new_n564), .C2(new_n568), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1081), .A2(new_n1089), .A3(new_n1083), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1034), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n996), .B2(G1996), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n555), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(new_n555), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1093), .A2(new_n1094), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1084), .A2(KEYINPUT122), .A3(new_n1090), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT122), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT61), .B(new_n1092), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1348), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1034), .A2(G2067), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT121), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1111), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1113), .B(new_n1114), .C1(new_n1010), .C2(G1348), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT60), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1112), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n608), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1119), .B2(new_n608), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n608), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1117), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(new_n1120), .A3(new_n608), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1109), .A2(new_n1123), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n608), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1116), .A2(new_n1130), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1092), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1079), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1023), .A2(new_n1020), .A3(G286), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1076), .A2(new_n1071), .A3(new_n1077), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1075), .A2(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1064), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1066), .A2(new_n1139), .A3(KEYINPUT63), .A4(new_n1134), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1076), .A2(new_n1049), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n719), .A2(new_n1044), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1039), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1035), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1030), .A2(new_n1149), .A3(new_n1032), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1025), .B(G8), .C1(new_n1029), .C2(G286), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1029), .A2(new_n1026), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1032), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1011), .A2(G171), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1141), .B(new_n1147), .C1(new_n1148), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n989), .B1(new_n1133), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n975), .A2(G1996), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT46), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n978), .A2(new_n982), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT47), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n975), .A2(G1986), .A3(G290), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT48), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1166), .A2(new_n1167), .B1(new_n986), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n980), .A2(new_n983), .A3(new_n704), .A4(new_n701), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(G2067), .B2(new_n759), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1172), .A2(new_n977), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1158), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g750(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n881), .A2(new_n693), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n954), .A2(new_n959), .ZN(new_n1179));
  NOR2_X1   g753(.A1(new_n1178), .A2(new_n1179), .ZN(G308));
  OR2_X1    g754(.A1(new_n1178), .A2(new_n1179), .ZN(G225));
endmodule


