//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(KEYINPUT3), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND3_X1  g051(.A1(new_n461), .A2(G2105), .A3(new_n465), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n462), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(G136), .B2(new_n467), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n477), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n469), .A2(new_n462), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n491), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n466), .B2(new_n492), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(KEYINPUT71), .B(KEYINPUT4), .C1(new_n466), .C2(new_n492), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n502), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT72), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n499), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n500), .B2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n502), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n511), .A2(KEYINPUT73), .A3(new_n501), .A4(new_n499), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT74), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n501), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n502), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(G651), .B1(G50), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n507), .A2(G89), .A3(new_n512), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(KEYINPUT75), .A3(new_n521), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n527), .A2(new_n531), .A3(G51), .A4(G543), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n511), .A2(new_n501), .A3(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n526), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(G168));
  AND2_X1   g114(.A1(new_n511), .A2(new_n501), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n507), .A2(G90), .A3(new_n512), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n527), .A2(new_n531), .A3(G543), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT76), .B(G52), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n544), .A2(KEYINPUT77), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT77), .B1(new_n544), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n543), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n540), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n542), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  INV_X1    g129(.A(new_n545), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n513), .A2(G81), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n545), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n517), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n513), .A2(G91), .B1(G651), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n550), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT78), .B(new_n543), .C1(new_n548), .C2(new_n549), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G301));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n526), .A2(new_n537), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n526), .B2(new_n537), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(G286));
  OAI21_X1  g154(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n545), .A2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n507), .A2(new_n512), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n513), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT81), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n540), .A2(new_n587), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n517), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G48), .B2(new_n522), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n513), .A2(new_n594), .A3(G86), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n586), .A2(new_n593), .A3(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n517), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G47), .B2(new_n545), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n582), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n513), .A2(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n540), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n542), .B1(new_n608), .B2(KEYINPUT83), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n555), .A2(KEYINPUT82), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n555), .B2(KEYINPUT82), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n604), .B1(new_n618), .B2(new_n603), .ZN(G284));
  AOI21_X1  g194(.A(new_n604), .B1(new_n618), .B2(new_n603), .ZN(G321));
  NOR2_X1   g195(.A1(G286), .A2(new_n603), .ZN(new_n621));
  XNOR2_X1  g196(.A(G299), .B(KEYINPUT85), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n603), .ZN(G297));
  AOI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n603), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  INV_X1    g201(.A(new_n558), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n603), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n617), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g206(.A1(new_n491), .A2(new_n472), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n467), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n478), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n462), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(G14), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(KEYINPUT17), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(new_n665), .B2(new_n661), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT87), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  OR2_X1    g244(.A1(new_n660), .A2(new_n661), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n669), .C1(new_n665), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(new_n683), .B(new_n682), .S(new_n675), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1981), .ZN(new_n686));
  INV_X1    g261(.A(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n690), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n690), .B2(new_n691), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(G229));
  XOR2_X1   g273(.A(KEYINPUT31), .B(G11), .Z(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT30), .B(G28), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n640), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n704));
  INV_X1    g279(.A(G34), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n705), .B2(new_n704), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n475), .B2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G2084), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(G32), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n478), .A2(G129), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n473), .A2(G105), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT98), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n467), .A2(G141), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT99), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT26), .ZN(new_n719));
  AND4_X1   g294(.A1(new_n712), .A2(new_n715), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n711), .B1(new_n720), .B2(new_n700), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  AOI211_X1 g297(.A(new_n703), .B(new_n710), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G162), .A2(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G29), .B2(G35), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT29), .B(G2090), .Z(new_n726));
  OAI221_X1 g301(.A(new_n723), .B1(new_n721), .B2(new_n722), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT25), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(new_n462), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n729), .B(new_n731), .C1(G139), .C2(new_n467), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G29), .B2(G33), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n709), .B2(new_n708), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n735), .B2(new_n734), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n558), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G16), .B2(G19), .ZN(new_n740));
  INV_X1    g315(.A(G1341), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n700), .A2(G27), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT100), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n494), .A2(new_n495), .ZN(new_n747));
  INV_X1    g322(.A(new_n493), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n747), .A2(new_n497), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n490), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n746), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT101), .Z(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G20), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G299), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n756), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n727), .A2(new_n744), .A3(new_n755), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n753), .A2(new_n754), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n617), .B2(new_n756), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1348), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n725), .A2(new_n726), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n700), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT96), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n478), .A2(G128), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT95), .Z(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(G116), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n467), .B2(G140), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2067), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n756), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n756), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n768), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G171), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G5), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n785), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n762), .A2(new_n763), .A3(new_n767), .A4(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G6), .B(G305), .S(G16), .Z(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT32), .B(G1981), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n756), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n756), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n756), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n756), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n795), .A2(new_n796), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT93), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NOR2_X1   g384(.A1(G25), .A2(G29), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n467), .A2(G131), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n478), .A2(G119), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(G29), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT90), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n756), .A2(G24), .ZN(new_n821));
  INV_X1    g396(.A(G290), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n756), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT91), .Z(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n825), .B2(G1986), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G1986), .B2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n809), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n792), .B1(new_n829), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(G311), .ZN(G150));
  INV_X1    g407(.A(KEYINPUT103), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n540), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(new_n542), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n507), .A2(G93), .A3(new_n512), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n545), .A2(G55), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n836), .A2(KEYINPUT102), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT102), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n627), .A2(new_n833), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n833), .ZN(new_n842));
  OAI211_X1 g417(.A(KEYINPUT103), .B(new_n835), .C1(new_n838), .C2(new_n839), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n558), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT38), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n618), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n840), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n720), .B(new_n751), .ZN(new_n856));
  INV_X1    g431(.A(new_n778), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(new_n857), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n855), .B(new_n732), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n732), .A2(new_n855), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n732), .A2(new_n855), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n862), .A2(new_n858), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n478), .A2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n462), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n467), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n633), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n816), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n861), .A2(new_n865), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n861), .B2(new_n865), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G160), .B(new_n640), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n873), .B2(new_n874), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n615), .B(new_n759), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n845), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n629), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n845), .B1(new_n617), .B2(G559), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n615), .B(G299), .ZN(new_n893));
  OAI211_X1 g468(.A(KEYINPUT105), .B(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(G288), .B(KEYINPUT106), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G305), .ZN(new_n897));
  XNOR2_X1  g472(.A(G303), .B(G290), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n891), .A2(new_n894), .A3(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n840), .A2(new_n603), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n883), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n603), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(new_n906), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(KEYINPUT107), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(G295));
  OR3_X1    g486(.A1(new_n908), .A2(KEYINPUT108), .A3(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G331));
  NAND2_X1  g489(.A1(new_n538), .A2(KEYINPUT79), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n526), .A2(new_n537), .A3(new_n576), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n550), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n544), .A2(new_n547), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT77), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n544), .A2(KEYINPUT77), .A3(new_n547), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  NAND4_X1  g499(.A1(G286), .A2(new_n923), .A3(new_n924), .A4(new_n543), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n572), .A2(G168), .A3(new_n573), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(KEYINPUT110), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT110), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n887), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n927), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n845), .A3(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n935), .A3(new_n884), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n845), .B1(new_n934), .B2(new_n928), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n934), .A2(KEYINPUT111), .A3(new_n845), .A4(new_n928), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n893), .B(new_n885), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n943), .B2(new_n899), .ZN(new_n944));
  INV_X1    g519(.A(new_n899), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n945), .B(new_n936), .C1(new_n941), .C2(new_n942), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT43), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n931), .A2(new_n884), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n939), .B2(new_n940), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n931), .B2(new_n935), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n899), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  AND4_X1   g527(.A1(KEYINPUT43), .A2(new_n951), .A3(new_n952), .A4(new_n946), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n943), .A2(new_n899), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n952), .A3(new_n946), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n946), .A3(new_n958), .A4(new_n952), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n954), .B1(new_n961), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g537(.A(G1384), .B1(new_n749), .B2(new_n750), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n475), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G164), .B2(G1384), .ZN(new_n970));
  INV_X1    g545(.A(new_n967), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT112), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n973), .A2(KEYINPUT114), .A3(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT114), .B1(new_n973), .B2(G1996), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n720), .ZN(new_n977));
  INV_X1    g552(.A(G2067), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n857), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n778), .A2(G2067), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(new_n720), .ZN(new_n983));
  INV_X1    g558(.A(new_n973), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n815), .B(new_n818), .Z(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT113), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n976), .B(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n981), .A2(new_n720), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n984), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n995), .B2(new_n998), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n816), .A2(new_n818), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n979), .B1(new_n986), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT126), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n984), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n963), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n967), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(G2084), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n751), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(new_n970), .A3(new_n967), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1011), .A2(KEYINPUT117), .B1(new_n783), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1010), .B2(G2084), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(G168), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1018), .A2(new_n1019), .A3(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n538), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(G8), .A3(new_n1018), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(KEYINPUT51), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n963), .B2(new_n967), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n801), .A2(G1976), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1026), .A2(KEYINPUT116), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1026), .A2(KEYINPUT115), .A3(new_n1027), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(KEYINPUT52), .A3(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n593), .A2(new_n585), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G1981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1026), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1034), .A2(new_n1039), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(G1971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1014), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1008), .A2(new_n1009), .A3(new_n1053), .A4(new_n967), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1025), .B(new_n1050), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1050), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(G8), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1048), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1013), .A2(new_n970), .A3(new_n754), .A4(new_n967), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1010), .A2(new_n788), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1060), .A2(KEYINPUT124), .A3(new_n1061), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT124), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1062), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n574), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1024), .A2(KEYINPUT62), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G286), .A2(new_n1025), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1021), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT118), .B(new_n1070), .C1(new_n1059), .C2(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1048), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1021), .A3(new_n1075), .A4(new_n1071), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1048), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1047), .A2(new_n1028), .A3(new_n801), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1040), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1078), .A2(new_n1055), .B1(new_n1080), .B2(new_n1026), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1069), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n967), .B1(new_n963), .B2(new_n1007), .ZN(new_n1084));
  NOR3_X1   g659(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT57), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1087), .A2(KEYINPUT57), .ZN(new_n1089));
  AND3_X1   g664(.A1(G299), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(G299), .B2(new_n1088), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1013), .A2(new_n970), .A3(new_n967), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1086), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n963), .A2(new_n967), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n963), .A2(KEYINPUT120), .A3(new_n967), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n978), .ZN(new_n1101));
  INV_X1    g676(.A(G1348), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1010), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n615), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1092), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1095), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1086), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1092), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1098), .A2(new_n1099), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1013), .A2(new_n970), .A3(new_n982), .A4(new_n967), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1115), .B1(new_n1120), .B2(new_n558), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n627), .B(new_n1114), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1109), .B(new_n1113), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT60), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1125));
  INV_X1    g700(.A(new_n615), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n615), .A4(new_n1103), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1106), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT123), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1065), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1060), .A2(KEYINPUT124), .A3(new_n1061), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1063), .B(KEYINPUT125), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n550), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n1066), .B2(new_n574), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1074), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n1136), .A3(G301), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT54), .B1(new_n1140), .B2(new_n1067), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1143), .B(new_n1106), .C1(new_n1123), .C2(new_n1129), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1131), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n1059), .A2(KEYINPUT62), .A3(new_n1067), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1024), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1082), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n990), .B1(G1986), .B2(G290), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n988), .B1(new_n973), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1006), .B1(new_n1149), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  INV_X1    g728(.A(G319), .ZN(new_n1155));
  NOR3_X1   g729(.A1(G401), .A2(new_n1155), .A3(G227), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n696), .A2(new_n697), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g731(.A(new_n1157), .B1(new_n878), .B2(new_n880), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n960), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n958), .B1(new_n944), .B2(new_n946), .ZN(new_n1160));
  INV_X1    g734(.A(new_n959), .ZN(new_n1161));
  OAI211_X1 g735(.A(new_n1158), .B(new_n1154), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g736(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g737(.A1(new_n1159), .A2(new_n1163), .ZN(G308));
  NAND2_X1  g738(.A1(new_n960), .A2(new_n1158), .ZN(G225));
endmodule


