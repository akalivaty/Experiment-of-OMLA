//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AND2_X1   g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n211), .A2(G20), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n209), .B(new_n213), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XOR2_X1   g0034(.A(G50), .B(G58), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(G45), .ZN(new_n241));
  NOR2_X1   g0041(.A1(new_n241), .A2(G1), .ZN(new_n242));
  AND2_X1   g0042(.A1(KEYINPUT5), .A2(G41), .ZN(new_n243));
  NOR2_X1   g0043(.A1(KEYINPUT5), .A2(G41), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n212), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(G257), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT5), .B(G41), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n249), .A2(new_n247), .A3(G274), .A4(new_n242), .ZN(new_n250));
  AND3_X1   g0050(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT80), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT80), .B1(new_n248), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(G33), .B2(G41), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(G250), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT79), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OAI211_X1 g0060(.A(G244), .B(new_n260), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G283), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n263), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n255), .B1(new_n259), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n253), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n253), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT6), .ZN(new_n278));
  INV_X1    g0078(.A(G97), .ZN(new_n279));
  INV_X1    g0079(.A(G107), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G97), .A2(G107), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(KEYINPUT6), .A3(G97), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n285), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n256), .A2(new_n257), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT7), .B1(new_n288), .B2(new_n204), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n267), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(G107), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n254), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT78), .B1(new_n298), .B2(new_n279), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT78), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n297), .A2(new_n300), .A3(G97), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n295), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n203), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI211_X1 g0105(.A(new_n299), .B(new_n301), .C1(new_n305), .C2(G97), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n275), .A2(new_n277), .A3(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n263), .A2(new_n269), .A3(new_n270), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT79), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n258), .B(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n247), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n248), .A2(new_n250), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT80), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n248), .A2(KEYINPUT80), .A3(new_n250), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(G200), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n253), .A2(new_n272), .A3(G190), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n318), .A2(new_n296), .A3(new_n306), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n297), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n305), .A2(new_n326), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n288), .A2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G68), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n265), .A2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G97), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT19), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT82), .ZN(new_n337));
  AND3_X1   g0137(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT19), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(new_n204), .ZN(new_n341));
  NOR3_X1   g0141(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n337), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n340), .B2(new_n204), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT82), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n336), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n295), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n328), .B(new_n329), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(G238), .B(new_n260), .C1(new_n256), .C2(new_n257), .ZN(new_n349));
  OAI211_X1 g0149(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n350));
  INV_X1    g0150(.A(G116), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n350), .C1(new_n265), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n255), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n203), .A2(G45), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT81), .A3(G250), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT81), .ZN(new_n356));
  AOI21_X1  g0156(.A(G274), .B1(new_n356), .B2(G250), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n247), .ZN(new_n359));
  AOI21_X1  g0159(.A(G169), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n359), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n360), .B1(new_n362), .B2(new_n276), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n348), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n330), .A2(G68), .B1(new_n334), .B2(new_n333), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n344), .A2(KEYINPUT82), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n337), .B(new_n342), .C1(new_n340), .C2(new_n204), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n327), .B1(new_n368), .B2(new_n295), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n353), .A2(G190), .A3(new_n359), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n353), .B2(new_n359), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G87), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n304), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n308), .A2(new_n320), .A3(new_n364), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n298), .A2(new_n280), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT25), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(G107), .B2(new_n305), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT84), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n204), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT22), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(KEYINPUT83), .A3(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n265), .A2(new_n351), .A3(G20), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT23), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n204), .B2(G107), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n280), .A2(KEYINPUT23), .A3(G20), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(KEYINPUT83), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT83), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n268), .A2(new_n394), .A3(new_n204), .A4(G87), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT22), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n383), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT24), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n347), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT22), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n386), .A2(new_n391), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT84), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n392), .A2(new_n383), .A3(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(KEYINPUT24), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT85), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT85), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n382), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n268), .A2(G250), .A3(new_n260), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G294), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n255), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n245), .A2(new_n247), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G264), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n417), .A3(new_n250), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n371), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT86), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(KEYINPUT86), .A3(new_n371), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n413), .A2(new_n255), .B1(new_n416), .B2(G264), .ZN(new_n423));
  INV_X1    g0223(.A(G190), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n250), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n378), .B1(new_n409), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT8), .B(G58), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n203), .B2(G20), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n302), .B1(new_n298), .B2(new_n429), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G68), .B1(new_n289), .B2(new_n291), .ZN(new_n433));
  INV_X1    g0233(.A(G58), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n217), .ZN(new_n435));
  NOR2_X1   g0235(.A1(G58), .A2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(G20), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n286), .A2(G159), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(KEYINPUT16), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n347), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n266), .A2(new_n204), .A3(new_n267), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT7), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n217), .B1(new_n446), .B2(new_n290), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n437), .A2(new_n438), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n432), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(G223), .B(new_n260), .C1(new_n256), .C2(new_n257), .ZN(new_n451));
  OAI211_X1 g0251(.A(G226), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n452));
  AND3_X1   g0252(.A1(KEYINPUT75), .A2(G33), .A3(G87), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT75), .B1(G33), .B2(G87), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n255), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n241), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n203), .A2(new_n459), .B1(new_n212), .B2(new_n246), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT64), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G45), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n463), .A3(new_n458), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n203), .A2(G274), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n460), .A2(G232), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n457), .A2(new_n276), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n465), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n247), .A2(G232), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n255), .B2(new_n456), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n467), .B1(new_n472), .B2(G169), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n428), .B1(new_n450), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n457), .A2(new_n276), .A3(new_n466), .ZN(new_n475));
  AOI21_X1  g0275(.A(G169), .B1(new_n457), .B2(new_n466), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n448), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n442), .B1(new_n433), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n295), .B1(new_n447), .B2(new_n439), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n431), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n481), .A3(KEYINPUT18), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT76), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n474), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n457), .A2(new_n424), .A3(new_n466), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n472), .B2(G200), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n450), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT17), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n441), .A2(new_n449), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n489), .A3(new_n431), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT77), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n477), .A2(new_n481), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT76), .A3(new_n428), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n484), .A2(new_n487), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n203), .A2(G20), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n324), .A2(G68), .A3(new_n347), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n332), .A2(KEYINPUT66), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT66), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n265), .B2(G20), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(G77), .A3(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n286), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n347), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n498), .B1(KEYINPUT11), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(KEYINPUT11), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n203), .A2(G13), .ZN(new_n507));
  NOR4_X1   g0307(.A1(new_n507), .A2(KEYINPUT12), .A3(new_n204), .A4(G68), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n321), .A2(new_n217), .A3(new_n323), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(KEYINPUT12), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n513));
  OAI211_X1 g0313(.A(G226), .B(new_n260), .C1(new_n256), .C2(new_n257), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n338), .A2(new_n339), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n255), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT13), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n460), .A2(G238), .B1(new_n464), .B2(new_n465), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n517), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g0321(.A(G169), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT13), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n522), .A2(KEYINPUT14), .B1(new_n526), .B2(new_n276), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT14), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n526), .B2(G169), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n512), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G200), .B1(new_n520), .B2(new_n521), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n524), .A2(G190), .A3(new_n525), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n511), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n496), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n499), .A2(new_n501), .ZN(new_n535));
  INV_X1    g0335(.A(new_n429), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n204), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(G150), .B2(new_n286), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n347), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n302), .A2(G50), .A3(new_n497), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(G50), .B2(new_n297), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT69), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT70), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n550), .A2(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(KEYINPUT9), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(new_n549), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n544), .A2(KEYINPUT69), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n550), .B(KEYINPUT9), .C1(new_n554), .C2(new_n548), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n460), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n468), .B1(new_n557), .B2(new_n216), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n268), .A2(G222), .A3(new_n260), .ZN(new_n559));
  INV_X1    g0359(.A(G77), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n268), .A2(G1698), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT65), .B(G223), .ZN(new_n562));
  OAI221_X1 g0362(.A(new_n559), .B1(new_n560), .B2(new_n268), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n558), .B1(new_n563), .B2(new_n255), .ZN(new_n564));
  OR3_X1    g0364(.A1(new_n564), .A2(KEYINPUT71), .A3(new_n371), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT71), .B1(new_n564), .B2(new_n371), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT10), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(G190), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n371), .B2(new_n564), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n553), .B2(new_n555), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n556), .A2(new_n569), .B1(new_n571), .B2(new_n567), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n564), .A2(new_n276), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n545), .C1(G169), .C2(new_n564), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n324), .A2(G77), .A3(new_n347), .A4(new_n497), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n326), .A2(new_n332), .B1(G20), .B2(G77), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n536), .A2(new_n286), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI221_X1 g0379(.A(new_n576), .B1(G77), .B2(new_n324), .C1(new_n579), .C2(new_n347), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n268), .A2(G232), .A3(new_n260), .ZN(new_n581));
  OAI221_X1 g0381(.A(new_n581), .B1(new_n280), .B2(new_n268), .C1(new_n561), .C2(new_n218), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n255), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n460), .A2(G244), .B1(new_n464), .B2(new_n465), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n371), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT68), .ZN(new_n586));
  OR3_X1    g0386(.A1(new_n580), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n580), .B2(new_n585), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n583), .A2(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G190), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n276), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n580), .C1(G169), .C2(new_n589), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n572), .A2(new_n575), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT72), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT72), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n572), .A2(new_n597), .A3(new_n575), .A4(new_n594), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n534), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n399), .A2(new_n407), .A3(new_n404), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n407), .B1(new_n399), .B2(new_n404), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n381), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n418), .A2(G179), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n274), .B2(new_n418), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n270), .B(new_n204), .C1(G33), .C2(new_n279), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n295), .C1(new_n204), .C2(G116), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n324), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n351), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n324), .A2(G116), .A3(new_n347), .A4(new_n303), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n268), .A2(G257), .A3(new_n260), .ZN(new_n615));
  INV_X1    g0415(.A(G303), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n268), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n255), .ZN(new_n618));
  INV_X1    g0418(.A(G270), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n250), .B1(new_n415), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n613), .A2(G169), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n613), .A2(KEYINPUT21), .A3(G169), .A4(new_n622), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n620), .B1(new_n255), .B2(new_n617), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n613), .A2(G179), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n613), .B1(G200), .B2(new_n622), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n424), .B2(new_n622), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n427), .A2(new_n599), .A3(new_n605), .A4(new_n632), .ZN(G372));
  INV_X1    g0433(.A(new_n572), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n474), .A2(new_n482), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n533), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n530), .B1(new_n593), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n492), .A2(new_n487), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n575), .B1(new_n634), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n605), .A2(new_n629), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n427), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n364), .A2(new_n377), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n308), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n327), .B(new_n375), .C1(new_n368), .C2(new_n295), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n373), .B1(new_n348), .B2(new_n363), .ZN(new_n648));
  INV_X1    g0448(.A(new_n308), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT26), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n646), .A2(new_n650), .B1(new_n348), .B2(new_n363), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n641), .B1(new_n599), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT87), .Z(G369));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n507), .A2(KEYINPUT27), .A3(G20), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT27), .B1(new_n507), .B2(G20), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n613), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n629), .A2(new_n631), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n613), .A3(new_n660), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT88), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(new_n667), .A3(new_n664), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n655), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n604), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n409), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n381), .B(new_n426), .C1(new_n600), .C2(new_n601), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n602), .A2(new_n660), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n605), .A2(new_n660), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n672), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n605), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n629), .A2(new_n660), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  NAND2_X1  g0482(.A1(new_n207), .A2(new_n458), .ZN(new_n683));
  INV_X1    g0483(.A(new_n342), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n210), .B2(new_n683), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n362), .A2(new_n627), .A3(G179), .A4(new_n423), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n273), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT30), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n689), .B2(new_n273), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n362), .A2(new_n627), .A3(G179), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n418), .A3(new_n273), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT31), .B1(new_n696), .B2(new_n660), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n695), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT89), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(KEYINPUT30), .B2(new_n690), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n693), .A2(new_n695), .A3(KEYINPUT89), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n660), .A2(KEYINPUT31), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT90), .B(new_n698), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n697), .ZN(new_n708));
  INV_X1    g0508(.A(new_n660), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n427), .A2(new_n605), .A3(new_n632), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n652), .A2(new_n713), .A3(new_n709), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n663), .B1(new_n602), .B2(new_n604), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n308), .A2(new_n320), .A3(new_n377), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n672), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n660), .B1(new_n718), .B2(new_n651), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n714), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n688), .B1(new_n721), .B2(G1), .ZN(G364));
  INV_X1    g0522(.A(new_n669), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n666), .A2(new_n655), .A3(new_n668), .ZN(new_n724));
  INV_X1    g0524(.A(new_n683), .ZN(new_n725));
  INV_X1    g0525(.A(G13), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n203), .B1(new_n727), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n725), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n207), .A2(new_n268), .ZN(new_n732));
  INV_X1    g0532(.A(G355), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(G116), .B2(new_n207), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n236), .A2(G45), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n207), .A2(new_n288), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n461), .A2(new_n463), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n211), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n734), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n254), .B1(G20), .B2(new_n274), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n731), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n424), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n276), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n279), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n204), .A2(new_n276), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n371), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n288), .B(new_n751), .C1(G68), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n424), .A2(new_n371), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n204), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n374), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n752), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n758), .A2(new_n753), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n560), .B1(new_n763), .B2(new_n280), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n752), .A2(new_n757), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n760), .B(new_n764), .C1(G50), .C2(new_n766), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n752), .A2(KEYINPUT91), .A3(new_n747), .ZN(new_n768));
  AOI21_X1  g0568(.A(KEYINPUT91), .B1(new_n752), .B2(new_n747), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G58), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n761), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n756), .A2(new_n767), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n763), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G329), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n759), .A2(new_n616), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(G326), .C2(new_n766), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n288), .B1(new_n762), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G294), .B2(new_n749), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT92), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT92), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(new_n755), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n771), .A2(G322), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n782), .A2(new_n785), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n777), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n746), .B1(new_n792), .B2(new_n743), .ZN(new_n793));
  INV_X1    g0593(.A(new_n742), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n665), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n730), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  INV_X1    g0597(.A(new_n712), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n594), .A2(new_n709), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n652), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n660), .B1(new_n643), .B2(new_n651), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n593), .A2(new_n660), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n580), .A2(new_n660), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n591), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(new_n805), .B2(new_n593), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n801), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n731), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n798), .B2(new_n807), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n766), .B1(new_n755), .B2(G150), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n774), .B2(new_n762), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n771), .B2(G143), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n750), .A2(new_n434), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n268), .B1(new_n773), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n763), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G68), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n215), .B2(new_n759), .ZN(new_n819));
  NOR4_X1   g0619(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n762), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G116), .A2(new_n821), .B1(new_n755), .B2(G283), .ZN(new_n822));
  INV_X1    g0622(.A(G294), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n783), .B2(new_n773), .C1(new_n823), .C2(new_n770), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n288), .B1(new_n759), .B2(new_n280), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n765), .A2(new_n616), .B1(new_n763), .B2(new_n374), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n824), .A2(new_n751), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n743), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n743), .A2(new_n740), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n729), .B(new_n725), .C1(new_n560), .C2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n828), .B(new_n830), .C1(new_n806), .C2(new_n741), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n809), .A2(new_n831), .ZN(G384));
  OR2_X1    g0632(.A1(new_n285), .A2(KEYINPUT35), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n285), .A2(KEYINPUT35), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n254), .A2(new_n204), .A3(new_n351), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT93), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n840));
  OAI21_X1  g0640(.A(G77), .B1(new_n434), .B2(new_n217), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n841), .A2(new_n210), .B1(G50), .B2(new_n217), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G1), .A3(new_n726), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT94), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n839), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT95), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n720), .A2(new_n599), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT101), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n720), .A2(new_n849), .A3(new_n599), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n641), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n522), .A2(KEYINPUT14), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n526), .A2(new_n528), .A3(G169), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(new_n276), .C2(new_n526), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n512), .B(new_n660), .C1(new_n854), .C2(new_n637), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n512), .A2(new_n660), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n530), .A2(new_n533), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n803), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n801), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n658), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n481), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n493), .A2(new_n863), .A3(new_n490), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n864), .A2(KEYINPUT97), .A3(KEYINPUT37), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT97), .B1(new_n864), .B2(KEYINPUT37), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n493), .A2(new_n863), .A3(new_n490), .A4(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT96), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n863), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n867), .A2(new_n871), .B1(new_n495), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n870), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n865), .B2(new_n866), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n873), .A2(KEYINPUT98), .A3(KEYINPUT38), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT97), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n864), .A2(KEYINPUT97), .A3(KEYINPUT37), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n871), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n495), .A2(new_n872), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n875), .A2(new_n881), .A3(KEYINPUT38), .A4(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT98), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n875), .A2(new_n881), .A3(new_n882), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n876), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n861), .A2(new_n889), .B1(new_n636), .B2(new_n658), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n876), .A2(new_n885), .A3(KEYINPUT39), .A4(new_n888), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n854), .A2(new_n512), .A3(new_n709), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n877), .A2(KEYINPUT100), .A3(new_n869), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n864), .A2(new_n896), .A3(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n863), .B1(new_n639), .B2(new_n635), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n883), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n891), .A2(new_n893), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n890), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n851), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n806), .A2(new_n858), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n698), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(new_n710), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n889), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n710), .A2(new_n698), .A3(new_n908), .ZN(new_n915));
  INV_X1    g0715(.A(new_n907), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n901), .A2(new_n915), .A3(new_n916), .A4(KEYINPUT40), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n599), .A2(new_n915), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(G330), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n906), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n923), .A2(KEYINPUT103), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n906), .A2(new_n922), .B1(new_n203), .B2(new_n727), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n923), .A2(KEYINPUT103), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n846), .B1(new_n926), .B2(new_n927), .ZN(G367));
  NAND2_X1  g0728(.A1(new_n671), .A2(new_n709), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n679), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n680), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n308), .A2(new_n709), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n307), .A2(new_n660), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n308), .A2(new_n320), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT42), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n929), .B1(new_n674), .B2(new_n931), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n649), .A2(new_n709), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n648), .B1(new_n647), .B2(new_n709), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n364), .A2(new_n647), .A3(new_n709), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n945), .A2(KEYINPUT105), .A3(new_n949), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n948), .B(KEYINPUT43), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n945), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n677), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n938), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT106), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(KEYINPUT106), .A3(new_n958), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n683), .B(KEYINPUT41), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n676), .A2(new_n680), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n967), .A2(new_n932), .A3(new_n669), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n669), .B1(new_n967), .B2(new_n932), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n681), .B2(new_n938), .ZN(new_n972));
  INV_X1    g0772(.A(new_n938), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n941), .A2(KEYINPUT44), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n929), .B(new_n938), .C1(new_n674), .C2(new_n931), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n681), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n970), .B(new_n721), .C1(new_n957), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n980), .A3(KEYINPUT107), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT108), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n677), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT107), .B1(new_n975), .B2(new_n980), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT109), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT107), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n981), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n990), .A2(new_n991), .A3(new_n985), .A4(new_n983), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n982), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n721), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n966), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n729), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(KEYINPUT110), .B(new_n966), .C1(new_n993), .C2(new_n994), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n964), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n946), .A2(new_n947), .A3(new_n742), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n744), .B1(new_n207), .B2(new_n325), .C1(new_n232), .C2(new_n736), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n731), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n763), .A2(new_n560), .ZN(new_n1003));
  INV_X1    g0803(.A(G137), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n268), .B1(new_n773), .B2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G143), .C2(new_n766), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n749), .A2(G68), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n771), .A2(G150), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n215), .A2(new_n762), .B1(new_n754), .B2(new_n774), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n759), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(G58), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n288), .B1(new_n762), .B2(new_n778), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(G116), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT46), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n1015), .B2(new_n1014), .C1(new_n280), .C2(new_n750), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(KEYINPUT111), .B(G311), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n766), .A2(new_n1019), .B1(new_n755), .B2(G294), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n773), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G97), .A2(new_n817), .B1(new_n1021), .B2(G317), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(new_n770), .C2(new_n616), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1012), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1002), .B1(new_n1025), .B2(new_n743), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1000), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n999), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(G387));
  AOI22_X1  g0830(.A1(G77), .A2(new_n1010), .B1(new_n1021), .B2(G150), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n268), .C1(new_n279), .C2(new_n763), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT114), .Z(new_n1033));
  NOR2_X1   g0833(.A1(new_n765), .A2(new_n774), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT115), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n750), .A2(new_n325), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n762), .A2(new_n217), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n754), .A2(new_n429), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1033), .B(new_n1039), .C1(new_n215), .C2(new_n770), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n268), .B1(new_n1021), .B2(G326), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n750), .A2(new_n778), .B1(new_n759), .B2(new_n823), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT116), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G322), .A2(new_n766), .B1(new_n821), .B2(G303), .ZN(new_n1044));
  INV_X1    g0844(.A(G317), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n754), .B2(new_n1018), .C1(new_n770), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1041), .B1(new_n351), .B2(new_n763), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1040), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n743), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n732), .A2(new_n685), .B1(G107), .B2(new_n207), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n229), .A2(new_n737), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n685), .ZN(new_n1057));
  AOI211_X1 g0857(.A(G45), .B(new_n1057), .C1(G68), .C2(G77), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n429), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n736), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1055), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n744), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n731), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1054), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n930), .B2(new_n742), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n970), .B2(new_n729), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n970), .A2(new_n721), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(KEYINPUT117), .A3(new_n725), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n721), .B2(new_n970), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT117), .B1(new_n1072), .B2(new_n725), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1071), .B1(new_n1074), .B2(new_n1075), .ZN(G393));
  INV_X1    g0876(.A(new_n993), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n981), .B(new_n957), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n683), .B1(new_n1078), .B2(new_n1072), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n728), .B1(new_n1078), .B2(KEYINPUT118), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(KEYINPUT118), .B2(new_n1078), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n973), .A2(new_n742), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n750), .A2(new_n560), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n288), .B(new_n1084), .C1(G87), .C2(new_n817), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G50), .A2(new_n755), .B1(new_n1010), .B2(G68), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n821), .A2(new_n536), .B1(new_n1021), .B2(G143), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(G150), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n770), .A2(new_n774), .B1(new_n1089), .B2(new_n765), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT51), .Z(new_n1091));
  AOI22_X1  g0891(.A1(G303), .A2(new_n755), .B1(new_n1021), .B2(G322), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n778), .B2(new_n759), .C1(new_n823), .C2(new_n762), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n288), .B1(new_n763), .B2(new_n280), .C1(new_n750), .C2(new_n351), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n770), .A2(new_n783), .B1(new_n1045), .B2(new_n765), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1088), .A2(new_n1091), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n743), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n744), .B1(new_n279), .B2(new_n207), .C1(new_n239), .C2(new_n736), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1083), .A2(new_n731), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1080), .A2(new_n1082), .A3(new_n1102), .ZN(G390));
  AND3_X1   g0903(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT120), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT120), .B1(new_n855), .B2(new_n857), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n805), .A2(new_n593), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n715), .A2(new_n717), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n645), .A2(new_n644), .A3(new_n308), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT26), .B1(new_n648), .B2(new_n649), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n364), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n709), .B(new_n1107), .C1(new_n1108), .C2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n1112), .B2(new_n860), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n901), .A2(new_n892), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n891), .A2(new_n903), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n799), .B1(new_n643), .B2(new_n651), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n858), .B1(new_n1117), .B2(new_n803), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n892), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n915), .A2(G330), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n907), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT121), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT121), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n891), .A2(new_n903), .B1(new_n1118), .B2(new_n892), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1122), .C1(new_n1126), .C2(new_n1115), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n711), .A2(G330), .A3(new_n806), .A4(new_n858), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1124), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n806), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1106), .B1(new_n1121), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1112), .A2(new_n860), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n711), .A2(G330), .A3(new_n806), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1122), .B1(new_n1135), .B2(new_n859), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1117), .A2(new_n803), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n599), .A2(G330), .A3(new_n915), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n851), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n725), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT122), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1143), .B(new_n725), .C1(new_n1130), .C2(new_n1140), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1130), .A2(new_n1140), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1124), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n729), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n829), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n731), .B1(new_n536), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G283), .A2(new_n766), .B1(new_n755), .B2(G107), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n279), .B2(new_n762), .C1(new_n770), .C2(new_n351), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n288), .B1(new_n759), .B2(new_n374), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n818), .B1(new_n823), .B2(new_n773), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1152), .A2(new_n1084), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(KEYINPUT123), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(KEYINPUT123), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n759), .A2(new_n1089), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT53), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n288), .B(new_n1160), .C1(G125), .C2(new_n1021), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1158), .A2(new_n1159), .B1(new_n749), .B2(G159), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n771), .A2(G132), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n765), .A2(new_n1164), .B1(new_n754), .B2(new_n1004), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n762), .A2(new_n1166), .B1(new_n763), .B2(new_n215), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1156), .A2(new_n1157), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1150), .B1(new_n1170), .B2(new_n743), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1116), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n741), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1148), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1146), .A2(new_n1175), .ZN(G378));
  OAI21_X1  g0976(.A(new_n731), .B1(G50), .B2(new_n1149), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n288), .B2(new_n458), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n763), .A2(new_n434), .B1(new_n773), .B2(new_n778), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n458), .B(new_n288), .C1(new_n759), .C2(new_n560), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G68), .C2(new_n749), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n765), .A2(new_n351), .B1(new_n754), .B2(new_n279), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n326), .B2(new_n821), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n280), .C2(new_n770), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n762), .A2(new_n1004), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n815), .A2(new_n754), .B1(new_n759), .B2(new_n1166), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G125), .C2(new_n766), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n1089), .B2(new_n750), .C1(new_n1164), .C2(new_n770), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n817), .A2(G159), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n1021), .C2(G124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1177), .B1(new_n1197), .B2(new_n743), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n658), .B1(new_n547), .B2(new_n549), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n572), .A2(new_n575), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n572), .B2(new_n575), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1200), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1205), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n1203), .A3(new_n1199), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1198), .B1(new_n1209), .B2(new_n741), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1209), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n917), .A2(G330), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n914), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n912), .B1(new_n889), .B2(new_n910), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1216), .A2(new_n1213), .A3(new_n1209), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n905), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n914), .A2(new_n1214), .A3(new_n1212), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n890), .A2(new_n904), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1209), .B1(new_n1216), .B2(new_n1213), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1211), .B1(new_n1223), .B2(new_n729), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n641), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n850), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n849), .B1(new_n720), .B2(new_n599), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(new_n1139), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1147), .B2(new_n1138), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1218), .A2(KEYINPUT124), .A3(new_n1222), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n905), .B(new_n1231), .C1(new_n1215), .C2(new_n1217), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n725), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1228), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1223), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1224), .B1(new_n1234), .B2(new_n1237), .ZN(G375));
  NAND2_X1  g1038(.A1(new_n1138), .A2(new_n729), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1106), .A2(new_n740), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n279), .A2(new_n759), .B1(new_n754), .B2(new_n351), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1036), .A2(new_n268), .A3(new_n1241), .A4(new_n1003), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G294), .A2(new_n766), .B1(new_n821), .B2(G107), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n616), .B2(new_n773), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G283), .B2(new_n771), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G132), .A2(new_n766), .B1(new_n821), .B2(G150), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1164), .B2(new_n773), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G137), .B2(new_n771), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n268), .B1(new_n763), .B2(new_n434), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n774), .A2(new_n759), .B1(new_n754), .B2(new_n1166), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(G50), .C2(new_n749), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1242), .A2(new_n1245), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n743), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n731), .B1(G68), .B2(new_n1149), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT125), .Z(new_n1255));
  NAND2_X1  g1055(.A1(new_n1240), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1239), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1235), .A2(new_n1138), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1140), .A2(new_n966), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(G381));
  OAI211_X1 g1061(.A(new_n796), .B(new_n1071), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(G378), .A2(G384), .A3(G381), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n995), .A2(new_n996), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n728), .A3(new_n998), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n962), .A2(new_n963), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1028), .B(G390), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G375), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1263), .A2(new_n1267), .A3(new_n1268), .ZN(G407));
  AOI22_X1  g1069(.A1(new_n1141), .A2(KEYINPUT122), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1174), .B1(new_n1270), .B2(new_n1144), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n659), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G407), .A2(G213), .A3(new_n1272), .ZN(G409));
  NAND3_X1  g1073(.A1(new_n1236), .A2(new_n966), .A3(new_n1223), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1230), .A2(new_n729), .A3(new_n1232), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1210), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1146), .A3(new_n1175), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(G375), .B2(new_n1271), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n659), .A2(G213), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1140), .A2(new_n725), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1138), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1228), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1228), .A3(new_n1281), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1280), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n809), .B(new_n831), .C1(new_n1286), .C2(new_n1257), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1285), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(new_n1283), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G384), .B(new_n1258), .C1(new_n1289), .C2(new_n1280), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1278), .A2(new_n1279), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1279), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(G2897), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1287), .A2(new_n1290), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1279), .A4(new_n1291), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1294), .A2(new_n1301), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G390), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1027), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT126), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G393), .A2(G396), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1262), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1309), .A2(new_n1308), .A3(new_n1262), .ZN(new_n1311));
  OAI22_X1  g1111(.A1(new_n1307), .A2(new_n1267), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(G390), .B1(new_n999), .B2(new_n1028), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1306), .A2(new_n1027), .A3(new_n1305), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1311), .A2(new_n1310), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1304), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G378), .B(new_n1224), .C1(new_n1237), .C2(new_n1234), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1296), .B1(new_n1322), .B2(new_n1277), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT62), .B1(new_n1323), .B2(new_n1291), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT62), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1292), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1320), .B(new_n1321), .C1(new_n1324), .C2(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1318), .A2(new_n1319), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1319), .B1(new_n1318), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1271), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1322), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1320), .B(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1291), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1291), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1317), .A2(new_n1332), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1320), .B1(new_n1322), .B2(new_n1331), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1338), .ZN(G402));
endmodule


