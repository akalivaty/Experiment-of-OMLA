

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733;

  AND2_X1 U372 ( .A1(n544), .A2(n543), .ZN(n569) );
  NOR2_X1 U373 ( .A1(n650), .A2(n653), .ZN(n520) );
  AND2_X1 U374 ( .A1(n661), .A2(n662), .ZN(n658) );
  XNOR2_X1 U375 ( .A(n581), .B(n519), .ZN(n648) );
  AND2_X1 U376 ( .A1(n536), .A2(n647), .ZN(n537) );
  NOR2_X1 U377 ( .A1(G902), .A2(n703), .ZN(n410) );
  XNOR2_X1 U378 ( .A(n714), .B(n371), .ZN(n350) );
  BUF_X1 U379 ( .A(G116), .Z(n351) );
  XNOR2_X1 U380 ( .A(n362), .B(KEYINPUT3), .ZN(n364) );
  XNOR2_X1 U381 ( .A(n350), .B(n420), .ZN(n606) );
  AND2_X4 U382 ( .A1(n597), .A2(n686), .ZN(n702) );
  XNOR2_X2 U383 ( .A(n462), .B(n360), .ZN(n721) );
  XNOR2_X2 U384 ( .A(n721), .B(n711), .ZN(n429) );
  XNOR2_X1 U385 ( .A(n439), .B(n438), .ZN(n680) );
  INV_X1 U386 ( .A(G953), .ZN(n725) );
  NOR2_X1 U387 ( .A1(n733), .A2(n732), .ZN(n547) );
  XNOR2_X2 U388 ( .A(n476), .B(KEYINPUT35), .ZN(n617) );
  NAND2_X1 U389 ( .A1(n558), .A2(n659), .ZN(n614) );
  NOR2_X1 U390 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U391 ( .A(n598), .B(n359), .ZN(n599) );
  NAND2_X2 U392 ( .A1(n518), .A2(n647), .ZN(n555) );
  INV_X1 U393 ( .A(n724), .ZN(n352) );
  INV_X1 U394 ( .A(n352), .ZN(n353) );
  INV_X1 U395 ( .A(KEYINPUT80), .ZN(n516) );
  INV_X1 U396 ( .A(KEYINPUT4), .ZN(n360) );
  XNOR2_X1 U397 ( .A(n457), .B(G475), .ZN(n458) );
  XNOR2_X1 U398 ( .A(n401), .B(n415), .ZN(n402) );
  XNOR2_X1 U399 ( .A(G113), .B(KEYINPUT11), .ZN(n444) );
  XNOR2_X1 U400 ( .A(G146), .B(G125), .ZN(n392) );
  XNOR2_X1 U401 ( .A(n545), .B(n357), .ZN(n584) );
  AND2_X1 U402 ( .A1(n601), .A2(G953), .ZN(n706) );
  XNOR2_X1 U403 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n534) );
  AND2_X1 U404 ( .A1(n675), .A2(n674), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n535), .B(n534), .ZN(n733) );
  NOR2_X1 U406 ( .A1(n678), .A2(n386), .ZN(n355) );
  AND2_X2 U407 ( .A1(n586), .A2(n356), .ZN(n724) );
  XNOR2_X2 U408 ( .A(n546), .B(KEYINPUT40), .ZN(n732) );
  AND2_X2 U409 ( .A1(n584), .A2(n639), .ZN(n546) );
  XNOR2_X1 U410 ( .A(n441), .B(n440), .ZN(n475) );
  NAND2_X1 U411 ( .A1(n500), .A2(n680), .ZN(n441) );
  XNOR2_X2 U412 ( .A(n484), .B(KEYINPUT32), .ZN(n611) );
  OR2_X2 U413 ( .A1(n510), .A2(n483), .ZN(n484) );
  XNOR2_X2 U414 ( .A(n668), .B(KEYINPUT6), .ZN(n548) );
  NOR2_X1 U415 ( .A1(n612), .A2(n585), .ZN(n356) );
  XOR2_X1 U416 ( .A(KEYINPUT69), .B(KEYINPUT39), .Z(n357) );
  XOR2_X1 U417 ( .A(KEYINPUT89), .B(KEYINPUT25), .Z(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT59), .B(KEYINPUT83), .ZN(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n395) );
  XNOR2_X1 U420 ( .A(n720), .B(n444), .ZN(n445) );
  XNOR2_X1 U421 ( .A(KEYINPUT75), .B(n724), .ZN(n587) );
  INV_X1 U422 ( .A(n646), .ZN(n585) );
  XNOR2_X1 U423 ( .A(KEYINPUT65), .B(G131), .ZN(n450) );
  XNOR2_X1 U424 ( .A(n456), .B(n455), .ZN(n598) );
  XNOR2_X1 U425 ( .A(n408), .B(n358), .ZN(n409) );
  BUF_X1 U426 ( .A(n618), .Z(n619) );
  OR2_X1 U427 ( .A1(n694), .A2(G902), .ZN(n422) );
  NAND2_X1 U428 ( .A1(n702), .A2(G475), .ZN(n600) );
  XNOR2_X1 U429 ( .A(n600), .B(n599), .ZN(n602) );
  XNOR2_X2 U430 ( .A(G143), .B(G128), .ZN(n462) );
  INV_X1 U431 ( .A(G101), .ZN(n711) );
  XOR2_X1 U432 ( .A(G110), .B(G107), .Z(n361) );
  XNOR2_X1 U433 ( .A(n361), .B(KEYINPUT74), .ZN(n712) );
  XNOR2_X1 U434 ( .A(n429), .B(n712), .ZN(n420) );
  XNOR2_X2 U435 ( .A(G119), .B(G116), .ZN(n362) );
  XNOR2_X1 U436 ( .A(G113), .B(KEYINPUT67), .ZN(n363) );
  XNOR2_X2 U437 ( .A(n364), .B(n363), .ZN(n430) );
  XNOR2_X1 U438 ( .A(G122), .B(G104), .ZN(n448) );
  XNOR2_X1 U439 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n365) );
  XNOR2_X1 U440 ( .A(n448), .B(n365), .ZN(n366) );
  XNOR2_X2 U441 ( .A(n430), .B(n366), .ZN(n714) );
  XNOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n367) );
  XNOR2_X1 U443 ( .A(n392), .B(n367), .ZN(n370) );
  NAND2_X1 U444 ( .A1(n725), .A2(G224), .ZN(n368) );
  XNOR2_X1 U445 ( .A(n368), .B(KEYINPUT77), .ZN(n369) );
  XNOR2_X1 U446 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U447 ( .A(G902), .B(KEYINPUT15), .ZN(n406) );
  INV_X1 U448 ( .A(n406), .ZN(n590) );
  OR2_X2 U449 ( .A1(n606), .A2(n590), .ZN(n378) );
  INV_X1 U450 ( .A(G902), .ZN(n434) );
  INV_X1 U451 ( .A(G237), .ZN(n373) );
  NAND2_X1 U452 ( .A1(n434), .A2(n373), .ZN(n379) );
  NAND2_X1 U453 ( .A1(n379), .A2(G210), .ZN(n376) );
  INV_X1 U454 ( .A(KEYINPUT78), .ZN(n374) );
  XNOR2_X1 U455 ( .A(n374), .B(KEYINPUT84), .ZN(n375) );
  XNOR2_X1 U456 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X2 U457 ( .A(n378), .B(n377), .ZN(n518) );
  NAND2_X1 U458 ( .A1(n379), .A2(G214), .ZN(n647) );
  INV_X1 U459 ( .A(KEYINPUT19), .ZN(n380) );
  XNOR2_X2 U460 ( .A(n555), .B(n380), .ZN(n561) );
  INV_X1 U461 ( .A(n561), .ZN(n387) );
  NAND2_X1 U462 ( .A1(G237), .A2(G234), .ZN(n382) );
  INV_X1 U463 ( .A(KEYINPUT14), .ZN(n381) );
  XNOR2_X1 U464 ( .A(n382), .B(n381), .ZN(n678) );
  NAND2_X1 U465 ( .A1(n725), .A2(G952), .ZN(n525) );
  INV_X1 U466 ( .A(G898), .ZN(n384) );
  NAND2_X1 U467 ( .A1(G953), .A2(G902), .ZN(n521) );
  INV_X1 U468 ( .A(n521), .ZN(n383) );
  NAND2_X1 U469 ( .A1(n384), .A2(n383), .ZN(n385) );
  AND2_X1 U470 ( .A1(n525), .A2(n385), .ZN(n386) );
  NAND2_X1 U471 ( .A1(n387), .A2(n355), .ZN(n389) );
  INV_X1 U472 ( .A(KEYINPUT0), .ZN(n388) );
  XNOR2_X1 U473 ( .A(n389), .B(n388), .ZN(n479) );
  INV_X1 U474 ( .A(n479), .ZN(n495) );
  XNOR2_X1 U475 ( .A(n495), .B(KEYINPUT85), .ZN(n500) );
  XOR2_X1 U476 ( .A(KEYINPUT64), .B(KEYINPUT8), .Z(n391) );
  NAND2_X1 U477 ( .A1(G234), .A2(n725), .ZN(n390) );
  XNOR2_X1 U478 ( .A(n391), .B(n390), .ZN(n468) );
  NAND2_X1 U479 ( .A1(G221), .A2(n468), .ZN(n405) );
  XNOR2_X1 U480 ( .A(n392), .B(KEYINPUT10), .ZN(n720) );
  XNOR2_X1 U481 ( .A(n720), .B(KEYINPUT68), .ZN(n403) );
  XOR2_X1 U482 ( .A(G110), .B(G137), .Z(n394) );
  XNOR2_X1 U483 ( .A(G128), .B(G119), .ZN(n393) );
  XNOR2_X1 U484 ( .A(n394), .B(n393), .ZN(n399) );
  INV_X1 U485 ( .A(n395), .ZN(n397) );
  XNOR2_X1 U486 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n396) );
  XNOR2_X1 U487 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U488 ( .A(n399), .B(n398), .ZN(n401) );
  INV_X1 U489 ( .A(KEYINPUT66), .ZN(n400) );
  XNOR2_X1 U490 ( .A(n400), .B(G140), .ZN(n415) );
  XNOR2_X1 U491 ( .A(n402), .B(n403), .ZN(n404) );
  XNOR2_X1 U492 ( .A(n405), .B(n404), .ZN(n703) );
  NAND2_X1 U493 ( .A1(n406), .A2(G234), .ZN(n407) );
  XNOR2_X1 U494 ( .A(n407), .B(KEYINPUT20), .ZN(n411) );
  NAND2_X1 U495 ( .A1(G217), .A2(n411), .ZN(n408) );
  XNOR2_X2 U496 ( .A(n410), .B(n409), .ZN(n661) );
  AND2_X1 U497 ( .A1(n411), .A2(G221), .ZN(n413) );
  XNOR2_X1 U498 ( .A(KEYINPUT90), .B(KEYINPUT21), .ZN(n412) );
  XNOR2_X1 U499 ( .A(n413), .B(n412), .ZN(n662) );
  XNOR2_X1 U500 ( .A(G137), .B(G134), .ZN(n414) );
  XNOR2_X1 U501 ( .A(n450), .B(n414), .ZN(n431) );
  XNOR2_X1 U502 ( .A(n431), .B(n415), .ZN(n723) );
  NAND2_X1 U503 ( .A1(n725), .A2(G227), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n416), .B(KEYINPUT86), .ZN(n418) );
  XNOR2_X1 U505 ( .A(G104), .B(G146), .ZN(n417) );
  XNOR2_X1 U506 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U507 ( .A(n723), .B(n419), .ZN(n421) );
  XNOR2_X1 U508 ( .A(n421), .B(n420), .ZN(n694) );
  XNOR2_X2 U509 ( .A(n422), .B(G469), .ZN(n531) );
  XNOR2_X2 U510 ( .A(n531), .B(KEYINPUT1), .ZN(n659) );
  NAND2_X1 U511 ( .A1(n658), .A2(n659), .ZN(n423) );
  XNOR2_X1 U512 ( .A(n423), .B(KEYINPUT107), .ZN(n437) );
  NOR2_X1 U513 ( .A1(G237), .A2(G953), .ZN(n424) );
  XNOR2_X1 U514 ( .A(n424), .B(KEYINPUT76), .ZN(n452) );
  NAND2_X1 U515 ( .A1(G210), .A2(n452), .ZN(n427) );
  XNOR2_X1 U516 ( .A(G146), .B(KEYINPUT5), .ZN(n425) );
  XNOR2_X1 U517 ( .A(n425), .B(KEYINPUT73), .ZN(n426) );
  XNOR2_X1 U518 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U519 ( .A(n429), .B(n428), .ZN(n433) );
  XNOR2_X1 U520 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U521 ( .A(n433), .B(n432), .ZN(n618) );
  NAND2_X1 U522 ( .A1(n618), .A2(n434), .ZN(n436) );
  XOR2_X1 U523 ( .A(G472), .B(KEYINPUT70), .Z(n435) );
  XNOR2_X2 U524 ( .A(n436), .B(n435), .ZN(n486) );
  BUF_X2 U525 ( .A(n486), .Z(n668) );
  NAND2_X1 U526 ( .A1(n437), .A2(n548), .ZN(n439) );
  XNOR2_X1 U527 ( .A(KEYINPUT108), .B(KEYINPUT33), .ZN(n438) );
  INV_X1 U528 ( .A(KEYINPUT34), .ZN(n440) );
  XOR2_X1 U529 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n443) );
  XNOR2_X1 U530 ( .A(KEYINPUT12), .B(KEYINPUT94), .ZN(n442) );
  XNOR2_X1 U531 ( .A(n443), .B(n442), .ZN(n446) );
  XNOR2_X1 U532 ( .A(n446), .B(n445), .ZN(n456) );
  XOR2_X1 U533 ( .A(G140), .B(KEYINPUT93), .Z(n447) );
  XNOR2_X1 U534 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U535 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U536 ( .A(G143), .B(n451), .Z(n454) );
  AND2_X1 U537 ( .A1(G214), .A2(n452), .ZN(n453) );
  XNOR2_X1 U538 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U539 ( .A1(G902), .A2(n598), .ZN(n459) );
  XNOR2_X1 U540 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n457) );
  XNOR2_X1 U541 ( .A(n459), .B(n458), .ZN(n504) );
  INV_X1 U542 ( .A(n504), .ZN(n502) );
  XOR2_X1 U543 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n461) );
  XNOR2_X1 U544 ( .A(G107), .B(KEYINPUT98), .ZN(n460) );
  XNOR2_X1 U545 ( .A(n461), .B(n460), .ZN(n472) );
  XNOR2_X1 U546 ( .A(G122), .B(KEYINPUT100), .ZN(n463) );
  XNOR2_X1 U547 ( .A(n463), .B(n462), .ZN(n467) );
  XOR2_X1 U548 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n465) );
  XNOR2_X1 U549 ( .A(n351), .B(G134), .ZN(n464) );
  XNOR2_X1 U550 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U551 ( .A(n467), .B(n466), .ZN(n470) );
  NAND2_X1 U552 ( .A1(G217), .A2(n468), .ZN(n469) );
  XNOR2_X1 U553 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U554 ( .A(n472), .B(n471), .ZN(n698) );
  NOR2_X1 U555 ( .A1(n698), .A2(G902), .ZN(n473) );
  XNOR2_X1 U556 ( .A(n473), .B(G478), .ZN(n501) );
  INV_X1 U557 ( .A(n501), .ZN(n503) );
  NAND2_X1 U558 ( .A1(n502), .A2(n503), .ZN(n567) );
  INV_X1 U559 ( .A(n567), .ZN(n474) );
  NAND2_X1 U560 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U561 ( .A1(n504), .A2(n501), .ZN(n477) );
  XNOR2_X1 U562 ( .A(n477), .B(KEYINPUT104), .ZN(n650) );
  INV_X1 U563 ( .A(n662), .ZN(n478) );
  NOR2_X1 U564 ( .A1(n650), .A2(n478), .ZN(n480) );
  NAND2_X1 U565 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U566 ( .A(n481), .B(KEYINPUT22), .ZN(n510) );
  NOR2_X1 U567 ( .A1(n548), .A2(n661), .ZN(n482) );
  NAND2_X1 U568 ( .A1(n482), .A2(n659), .ZN(n483) );
  INV_X1 U569 ( .A(KEYINPUT106), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n486), .B(n485), .ZN(n536) );
  NOR2_X1 U571 ( .A1(n536), .A2(n661), .ZN(n487) );
  INV_X1 U572 ( .A(n659), .ZN(n507) );
  NAND2_X1 U573 ( .A1(n487), .A2(n507), .ZN(n488) );
  OR2_X1 U574 ( .A1(n510), .A2(n488), .ZN(n634) );
  NAND2_X1 U575 ( .A1(n611), .A2(n634), .ZN(n489) );
  NOR2_X2 U576 ( .A1(n617), .A2(n489), .ZN(n490) );
  XNOR2_X1 U577 ( .A(n490), .B(KEYINPUT44), .ZN(n514) );
  AND2_X1 U578 ( .A1(n658), .A2(n659), .ZN(n492) );
  INV_X1 U579 ( .A(n668), .ZN(n491) );
  NAND2_X1 U580 ( .A1(n492), .A2(n491), .ZN(n494) );
  INV_X1 U581 ( .A(KEYINPUT91), .ZN(n493) );
  XNOR2_X1 U582 ( .A(n494), .B(n493), .ZN(n670) );
  OR2_X1 U583 ( .A1(n495), .A2(n670), .ZN(n497) );
  XNOR2_X1 U584 ( .A(KEYINPUT92), .B(KEYINPUT31), .ZN(n496) );
  XNOR2_X1 U585 ( .A(n497), .B(n496), .ZN(n642) );
  NAND2_X1 U586 ( .A1(n658), .A2(n668), .ZN(n498) );
  INV_X1 U587 ( .A(n531), .ZN(n541) );
  NOR2_X1 U588 ( .A1(n498), .A2(n541), .ZN(n499) );
  AND2_X1 U589 ( .A1(n500), .A2(n499), .ZN(n630) );
  OR2_X1 U590 ( .A1(n642), .A2(n630), .ZN(n506) );
  NOR2_X1 U591 ( .A1(n502), .A2(n501), .ZN(n643) );
  XNOR2_X1 U592 ( .A(KEYINPUT102), .B(n643), .ZN(n583) );
  OR2_X1 U593 ( .A1(n504), .A2(n503), .ZN(n553) );
  INV_X1 U594 ( .A(n553), .ZN(n639) );
  NOR2_X1 U595 ( .A1(n583), .A2(n639), .ZN(n505) );
  XNOR2_X1 U596 ( .A(KEYINPUT103), .B(n505), .ZN(n563) );
  INV_X1 U597 ( .A(n563), .ZN(n652) );
  NAND2_X1 U598 ( .A1(n506), .A2(n563), .ZN(n511) );
  INV_X1 U599 ( .A(n661), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n548), .A2(n542), .ZN(n508) );
  NAND2_X1 U601 ( .A1(n508), .A2(n507), .ZN(n509) );
  OR2_X1 U602 ( .A1(n510), .A2(n509), .ZN(n626) );
  NAND2_X1 U603 ( .A1(n511), .A2(n626), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n512), .B(KEYINPUT105), .ZN(n513) );
  NAND2_X1 U605 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U606 ( .A(n515), .B(KEYINPUT45), .ZN(n594) );
  NAND2_X1 U607 ( .A1(n594), .A2(n590), .ZN(n517) );
  XNOR2_X1 U608 ( .A(n517), .B(n516), .ZN(n589) );
  BUF_X2 U609 ( .A(n518), .Z(n581) );
  INV_X1 U610 ( .A(KEYINPUT38), .ZN(n519) );
  NAND2_X1 U611 ( .A1(n648), .A2(n647), .ZN(n653) );
  XNOR2_X1 U612 ( .A(n520), .B(KEYINPUT41), .ZN(n672) );
  INV_X1 U613 ( .A(n672), .ZN(n533) );
  NOR2_X1 U614 ( .A1(n678), .A2(n521), .ZN(n522) );
  XNOR2_X1 U615 ( .A(n522), .B(KEYINPUT109), .ZN(n523) );
  NOR2_X1 U616 ( .A1(G900), .A2(n523), .ZN(n524) );
  XNOR2_X1 U617 ( .A(n524), .B(KEYINPUT110), .ZN(n527) );
  NOR2_X1 U618 ( .A1(n678), .A2(n525), .ZN(n526) );
  NOR2_X1 U619 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U620 ( .A(KEYINPUT79), .B(n528), .ZN(n529) );
  NAND2_X1 U621 ( .A1(n529), .A2(n662), .ZN(n539) );
  NOR2_X1 U622 ( .A1(n661), .A2(n539), .ZN(n549) );
  AND2_X1 U623 ( .A1(n536), .A2(n549), .ZN(n530) );
  XNOR2_X1 U624 ( .A(KEYINPUT28), .B(n530), .ZN(n532) );
  AND2_X1 U625 ( .A1(n532), .A2(n531), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n533), .A2(n560), .ZN(n535) );
  INV_X1 U627 ( .A(KEYINPUT30), .ZN(n538) );
  XNOR2_X1 U628 ( .A(n538), .B(n537), .ZN(n540) );
  NOR2_X1 U629 ( .A1(n540), .A2(n539), .ZN(n544) );
  NOR2_X1 U630 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U631 ( .A1(n569), .A2(n648), .ZN(n545) );
  XNOR2_X1 U632 ( .A(n547), .B(KEYINPUT46), .ZN(n559) );
  INV_X1 U633 ( .A(KEYINPUT111), .ZN(n551) );
  NAND2_X1 U634 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U635 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U636 ( .A(KEYINPUT112), .B(n554), .ZN(n579) );
  XOR2_X1 U637 ( .A(KEYINPUT114), .B(n579), .Z(n556) );
  NOR2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U639 ( .A(n557), .B(KEYINPUT36), .ZN(n558) );
  NAND2_X1 U640 ( .A1(n559), .A2(n614), .ZN(n575) );
  INV_X1 U641 ( .A(KEYINPUT72), .ZN(n570) );
  NOR2_X1 U642 ( .A1(n570), .A2(KEYINPUT47), .ZN(n565) );
  INV_X1 U643 ( .A(n560), .ZN(n562) );
  NOR2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n637) );
  NAND2_X1 U645 ( .A1(n563), .A2(n637), .ZN(n564) );
  XNOR2_X1 U646 ( .A(n565), .B(n564), .ZN(n573) );
  INV_X1 U647 ( .A(n581), .ZN(n566) );
  NOR2_X1 U648 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U649 ( .A1(n569), .A2(n568), .ZN(n616) );
  NAND2_X1 U650 ( .A1(n570), .A2(KEYINPUT47), .ZN(n571) );
  AND2_X1 U651 ( .A1(n616), .A2(n571), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X2 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U654 ( .A(n576), .B(KEYINPUT48), .ZN(n586) );
  INV_X1 U655 ( .A(n647), .ZN(n577) );
  NOR2_X1 U656 ( .A1(n659), .A2(n577), .ZN(n578) );
  NAND2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U658 ( .A(KEYINPUT43), .B(n580), .Z(n582) );
  NOR2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n612) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n646) );
  INV_X1 U661 ( .A(n587), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n590), .A2(KEYINPUT2), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n724), .A2(KEYINPUT2), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT81), .ZN(n596) );
  BUF_X1 U667 ( .A(n594), .Z(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n686) );
  INV_X1 U669 ( .A(G952), .ZN(n601) );
  NOR2_X2 U670 ( .A1(n602), .A2(n706), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U672 ( .A1(n702), .A2(G210), .ZN(n608) );
  XOR2_X1 U673 ( .A(KEYINPUT124), .B(KEYINPUT54), .Z(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(KEYINPUT55), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U676 ( .A(n608), .B(n607), .ZN(n609) );
  NOR2_X2 U677 ( .A1(n609), .A2(n706), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n610), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U679 ( .A(n611), .B(G119), .ZN(G21) );
  XOR2_X1 U680 ( .A(G140), .B(n612), .Z(G42) );
  XOR2_X1 U681 ( .A(G125), .B(KEYINPUT37), .Z(n613) );
  XNOR2_X1 U682 ( .A(n614), .B(n613), .ZN(G27) );
  XOR2_X1 U683 ( .A(G143), .B(KEYINPUT117), .Z(n615) );
  XNOR2_X1 U684 ( .A(n616), .B(n615), .ZN(G45) );
  XOR2_X1 U685 ( .A(n617), .B(G122), .Z(G24) );
  NAND2_X1 U686 ( .A1(n702), .A2(G472), .ZN(n621) );
  XOR2_X1 U687 ( .A(KEYINPUT62), .B(n619), .Z(n620) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X2 U689 ( .A1(n622), .A2(n706), .ZN(n625) );
  XNOR2_X1 U690 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(KEYINPUT82), .ZN(n624) );
  XNOR2_X1 U692 ( .A(n625), .B(n624), .ZN(G57) );
  INV_X1 U693 ( .A(n626), .ZN(n627) );
  XOR2_X1 U694 ( .A(G101), .B(n627), .Z(G3) );
  XNOR2_X1 U695 ( .A(G104), .B(KEYINPUT116), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n630), .A2(n639), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(G6) );
  XOR2_X1 U698 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U699 ( .A1(n630), .A2(n643), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U701 ( .A(G107), .B(n633), .ZN(G9) );
  XNOR2_X1 U702 ( .A(G110), .B(n634), .ZN(G12) );
  XOR2_X1 U703 ( .A(G128), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U704 ( .A1(n637), .A2(n643), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(G30) );
  NAND2_X1 U706 ( .A1(n637), .A2(n639), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n638), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n642), .A2(n639), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n640), .B(KEYINPUT118), .ZN(n641) );
  XNOR2_X1 U710 ( .A(G113), .B(n641), .ZN(G15) );
  XOR2_X1 U711 ( .A(n351), .B(KEYINPUT119), .Z(n645) );
  NAND2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n645), .B(n644), .ZN(G18) );
  XNOR2_X1 U714 ( .A(G134), .B(n646), .ZN(G36) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT121), .B(n651), .Z(n655) );
  NOR2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n657) );
  INV_X1 U720 ( .A(n680), .ZN(n656) );
  OR2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n675) );
  NOR2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U724 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(n663), .Z(n664) );
  XNOR2_X1 U726 ( .A(n664), .B(KEYINPUT120), .ZN(n665) );
  NOR2_X1 U727 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n671), .ZN(n673) );
  OR2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U732 ( .A(n354), .B(KEYINPUT52), .ZN(n676) );
  XNOR2_X1 U733 ( .A(KEYINPUT122), .B(n676), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U735 ( .A1(G952), .A2(n679), .ZN(n682) );
  NAND2_X1 U736 ( .A1(n533), .A2(n680), .ZN(n681) );
  NAND2_X1 U737 ( .A1(n682), .A2(n681), .ZN(n688) );
  NAND2_X1 U738 ( .A1(n353), .A2(n595), .ZN(n684) );
  INV_X1 U739 ( .A(KEYINPUT2), .ZN(n683) );
  NAND2_X1 U740 ( .A1(n684), .A2(n683), .ZN(n685) );
  AND2_X1 U741 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U742 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT123), .ZN(n690) );
  NOR2_X1 U744 ( .A1(G953), .A2(n690), .ZN(n691) );
  XNOR2_X1 U745 ( .A(KEYINPUT53), .B(n691), .ZN(G75) );
  NAND2_X1 U746 ( .A1(n702), .A2(G469), .ZN(n696) );
  XNOR2_X1 U747 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n692), .B(KEYINPUT57), .ZN(n693) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U751 ( .A1(n706), .A2(n697), .ZN(G54) );
  NAND2_X1 U752 ( .A1(n702), .A2(G478), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n698), .B(KEYINPUT126), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n706), .A2(n701), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n702), .A2(G217), .ZN(n704) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U759 ( .A1(n595), .A2(n725), .ZN(n710) );
  NAND2_X1 U760 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n708), .A2(G898), .ZN(n709) );
  NAND2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n718) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U766 ( .A1(G898), .A2(n725), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U769 ( .A(KEYINPUT127), .B(n719), .Z(G69) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n723), .B(n722), .ZN(n727) );
  XOR2_X1 U772 ( .A(n727), .B(n353), .Z(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(n725), .ZN(n731) );
  XNOR2_X1 U774 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U776 ( .A1(G953), .A2(n729), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U778 ( .A(n732), .B(G131), .Z(G33) );
  XOR2_X1 U779 ( .A(n733), .B(G137), .Z(G39) );
endmodule

