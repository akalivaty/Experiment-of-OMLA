//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G127gat), .A2(G134gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G127gat), .A2(G134gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n208), .B2(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G127gat), .A2(G134gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT66), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n217), .A2(new_n218), .A3(new_n206), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n217), .B2(new_n206), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT73), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n208), .A2(new_n207), .A3(new_n210), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT66), .B1(new_n214), .B2(new_n215), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n206), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n217), .A2(new_n218), .A3(new_n206), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT73), .A3(new_n209), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT2), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G155gat), .B(G162gat), .Z(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n238), .C1(new_n239), .C2(KEYINPUT72), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n233), .A3(new_n234), .ZN(new_n241));
  XNOR2_X1  g040(.A(G155gat), .B(G162gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n233), .A2(KEYINPUT72), .A3(new_n234), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT3), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n240), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n230), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n223), .A2(new_n230), .A3(new_n247), .A4(KEYINPUT74), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(new_n244), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n209), .C1(new_n219), .C2(new_n220), .ZN(new_n254));
  OR3_X1    g053(.A1(new_n254), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT76), .B1(new_n254), .B2(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n252), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n263));
  INV_X1    g062(.A(new_n253), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n223), .A2(new_n230), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n254), .ZN(new_n266));
  INV_X1    g065(.A(new_n261), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT77), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n229), .A2(new_n209), .A3(new_n253), .A4(new_n257), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n263), .A4(new_n261), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n270), .B1(new_n252), .B2(new_n275), .ZN(new_n276));
  AOI211_X1 g075(.A(KEYINPUT77), .B(new_n274), .C1(new_n250), .C2(new_n251), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G1gat), .B(G29gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G85gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n269), .B(new_n282), .C1(new_n276), .C2(new_n277), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n252), .A2(new_n275), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT77), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n252), .A2(new_n270), .A3(new_n275), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n291), .A2(new_n292), .B1(new_n262), .B2(new_n268), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n282), .B(KEYINPUT80), .Z(new_n294));
  OAI211_X1 g093(.A(new_n289), .B(new_n284), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n278), .A2(KEYINPUT83), .A3(new_n283), .A4(new_n285), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301));
  INV_X1    g100(.A(G211gat), .ZN(new_n302));
  INV_X1    g101(.A(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n300), .A3(new_n304), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n315));
  OAI22_X1  g114(.A1(new_n315), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n313), .B(new_n314), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  AND2_X1   g119(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n311), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n323), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n321), .ZN(new_n328));
  INV_X1    g127(.A(new_n314), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(KEYINPUT23), .B2(new_n312), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n331), .B(new_n332), .C1(G169gat), .C2(G176gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n328), .A2(KEYINPUT25), .A3(new_n330), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  NOR3_X1   g134(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(KEYINPUT65), .A3(new_n314), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n336), .A2(new_n340), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n342), .A2(KEYINPUT28), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT28), .B1(new_n342), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n339), .B(new_n341), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n335), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n335), .B2(new_n346), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n310), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n346), .A3(new_n347), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n308), .A2(new_n309), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n344), .A2(new_n345), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n339), .A2(new_n341), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(new_n325), .B2(new_n334), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n352), .B(new_n353), .C1(new_n356), .C2(new_n349), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(new_n357), .A3(KEYINPUT69), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n359), .B(new_n310), .C1(new_n348), .C2(new_n350), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT37), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n299), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n351), .A2(new_n357), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT38), .B1(new_n364), .B2(KEYINPUT37), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT38), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n358), .A2(KEYINPUT37), .A3(new_n360), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n299), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n358), .B2(new_n360), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n288), .A2(new_n295), .A3(new_n296), .A4(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n360), .A3(new_n370), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n299), .A2(KEYINPUT30), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n361), .A2(KEYINPUT70), .A3(new_n377), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n371), .A2(KEYINPUT30), .ZN(new_n383));
  INV_X1    g182(.A(new_n294), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n382), .A2(new_n383), .B1(new_n278), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT40), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT39), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n272), .A2(new_n273), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n252), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n267), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n265), .A2(new_n254), .A3(new_n261), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT82), .Z(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AOI211_X1 g192(.A(KEYINPUT39), .B(new_n261), .C1(new_n252), .C2(new_n388), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n394), .A2(KEYINPUT81), .A3(new_n384), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n387), .A3(new_n267), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(new_n294), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT81), .B1(new_n394), .B2(new_n384), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n396), .A3(new_n294), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n400), .A2(new_n401), .B1(new_n392), .B2(new_n390), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n385), .B(new_n399), .C1(new_n402), .C2(KEYINPUT40), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n353), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n253), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n310), .B1(new_n246), .B2(KEYINPUT29), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n253), .A2(new_n406), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n353), .B1(new_n412), .B2(new_n404), .ZN(new_n413));
  OAI21_X1  g212(.A(G22gat), .B1(new_n413), .B2(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n410), .B2(KEYINPUT79), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n417), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(new_n411), .A3(new_n414), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n418), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n373), .A2(new_n403), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n289), .A2(new_n284), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n293), .A2(new_n282), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n286), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT70), .B1(new_n361), .B2(new_n377), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n379), .B(new_n376), .C1(new_n358), .C2(new_n360), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n374), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT71), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT71), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n374), .C1(new_n431), .C2(new_n432), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n436), .A3(new_n383), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n426), .ZN(new_n440));
  XOR2_X1   g239(.A(G15gat), .B(G43gat), .Z(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G227gat), .ZN(new_n445));
  INV_X1    g244(.A(G233gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n335), .A2(new_n346), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n221), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n229), .A2(new_n209), .B1(new_n335), .B2(new_n346), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n221), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n229), .A2(new_n209), .A3(new_n335), .A4(new_n346), .ZN(new_n455));
  INV_X1    g254(.A(new_n447), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n455), .A3(new_n459), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n455), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT33), .B1(new_n463), .B2(new_n447), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n458), .B(new_n460), .C1(new_n464), .C2(new_n444), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT32), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT68), .B(KEYINPUT36), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n462), .A2(new_n465), .A3(new_n469), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n462), .B2(new_n465), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n439), .A2(new_n440), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n426), .A2(new_n468), .A3(new_n470), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n474), .A2(new_n475), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n426), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT35), .B1(new_n439), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n288), .A2(new_n295), .A3(new_n296), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n382), .A2(new_n383), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n486), .A2(new_n478), .A3(KEYINPUT35), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n427), .A2(new_n477), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(G1gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT16), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(G1gat), .B2(new_n490), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(G8gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT87), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  AND2_X1   g296(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G43gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT15), .B1(new_n504), .B2(G50gat), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n504), .B2(G50gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  OR3_X1    g307(.A1(new_n508), .A2(KEYINPUT86), .A3(G43gat), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n504), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT86), .B1(new_n508), .B2(G43gat), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT85), .B1(new_n504), .B2(G50gat), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n513), .A2(new_n514), .B1(new_n500), .B2(new_n502), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n507), .B1(new_n515), .B2(new_n506), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT17), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT88), .Z(new_n521));
  OR2_X1    g320(.A1(new_n495), .A2(new_n516), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n519), .A2(KEYINPUT18), .A3(new_n521), .A4(new_n522), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n495), .B(new_n516), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n521), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT12), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n525), .A2(new_n538), .A3(new_n526), .A4(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n489), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  OR2_X1    g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G57gat), .B(G64gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT91), .ZN(new_n549));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n545), .B1(new_n550), .B2(KEYINPUT90), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(KEYINPUT90), .B2(new_n550), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n544), .A2(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n495), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT95), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n558), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G127gat), .B(G155gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT94), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT93), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n565), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G183gat), .B(G211gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n563), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT96), .Z(new_n573));
  XOR2_X1   g372(.A(G134gat), .B(G162gat), .Z(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(G85gat), .A2(G92gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G99gat), .B(G106gat), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n580), .A3(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n578), .B1(new_n516), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT97), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n518), .A2(new_n517), .A3(new_n590), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n577), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n575), .B1(new_n594), .B2(KEYINPUT98), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n577), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n594), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(KEYINPUT98), .A3(new_n596), .A4(new_n575), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n571), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n589), .A2(KEYINPUT99), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n549), .A2(new_n554), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n590), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n608), .B1(new_n552), .B2(new_n553), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n590), .A3(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n555), .A2(new_n617), .A3(new_n590), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n604), .A2(new_n605), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n590), .B1(new_n609), .B2(new_n603), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n610), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(KEYINPUT100), .A3(new_n617), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n618), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n611), .B1(new_n626), .B2(KEYINPUT101), .ZN(new_n627));
  INV_X1    g426(.A(new_n618), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT100), .B1(new_n624), .B2(new_n617), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n622), .B(KEYINPUT10), .C1(new_n606), .C2(new_n610), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n613), .B(new_n616), .C1(new_n627), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n611), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n613), .ZN(new_n636));
  INV_X1    g435(.A(new_n616), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n602), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n542), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n430), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n491), .ZN(G1324gat));
  AND2_X1   g442(.A1(new_n542), .A2(new_n640), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n486), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n486), .ZN(new_n649));
  OAI21_X1  g448(.A(G8gat), .B1(new_n641), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT102), .B1(new_n648), .B2(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(G1325gat));
  AOI21_X1  g455(.A(G15gat), .B1(new_n644), .B2(new_n480), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n476), .A2(new_n472), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n476), .B2(new_n472), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G15gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT104), .Z(new_n664));
  AOI21_X1  g463(.A(new_n657), .B1(new_n644), .B2(new_n664), .ZN(G1326gat));
  NAND3_X1  g464(.A1(new_n542), .A2(new_n440), .A3(new_n640), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NOR3_X1   g467(.A1(new_n639), .A2(new_n571), .A3(new_n601), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n542), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n430), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n501), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n373), .A2(new_n403), .A3(new_n426), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n278), .A2(new_n283), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n284), .A3(new_n289), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n437), .B1(new_n676), .B2(new_n286), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n661), .B1(new_n677), .B2(new_n426), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT35), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n479), .A2(new_n482), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n485), .A2(new_n487), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n674), .A2(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n439), .A2(new_n440), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n427), .A2(new_n686), .A3(new_n661), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(KEYINPUT106), .C1(new_n681), .C2(new_n682), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n601), .A2(KEYINPUT44), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n489), .B2(new_n601), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n639), .ZN(new_n693));
  INV_X1    g492(.A(new_n571), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n540), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n430), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n698), .B2(KEYINPUT107), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n673), .B1(new_n699), .B2(new_n700), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n670), .A2(new_n497), .A3(new_n486), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT46), .Z(new_n703));
  OAI21_X1  g502(.A(G36gat), .B1(new_n697), .B2(new_n649), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n474), .A2(new_n475), .A3(G43gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n542), .A2(new_n669), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n696), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n690), .B2(new_n691), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n504), .B1(new_n712), .B2(new_n662), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n661), .B(new_n711), .C1(new_n690), .C2(new_n691), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(KEYINPUT108), .A3(new_n504), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n706), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  OAI21_X1  g518(.A(G43gat), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n697), .A2(KEYINPUT110), .A3(new_n661), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT47), .B(new_n710), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1330gat));
  AND4_X1   g522(.A1(new_n508), .A2(new_n542), .A3(new_n440), .A4(new_n669), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n712), .A2(new_n440), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(G50gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g526(.A1(new_n685), .A2(new_n688), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n693), .A2(new_n602), .A3(new_n540), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n430), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT111), .B(G57gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n649), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n730), .B2(new_n661), .ZN(new_n739));
  INV_X1    g538(.A(G71gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n480), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n730), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n730), .A2(new_n426), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT113), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n541), .B2(new_n694), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n540), .A2(new_n571), .A3(KEYINPUT114), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n693), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n692), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n430), .ZN(new_n754));
  INV_X1    g553(.A(new_n683), .ZN(new_n755));
  INV_X1    g554(.A(new_n601), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n749), .B2(new_n750), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT51), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n755), .B2(new_n757), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n693), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n582), .A3(new_n671), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n754), .A2(new_n763), .ZN(G1336gat));
  NOR2_X1   g563(.A1(new_n649), .A2(G92gat), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n753), .B2(new_n649), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n758), .A2(KEYINPUT115), .A3(new_n760), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n760), .B1(new_n758), .B2(KEYINPUT115), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n769), .A2(new_n639), .A3(new_n770), .A4(new_n765), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(G1337gat));
  AND2_X1   g573(.A1(new_n692), .A2(new_n752), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(G99gat), .A3(new_n662), .ZN(new_n776));
  AOI21_X1  g575(.A(G99gat), .B1(new_n762), .B2(new_n480), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(G1338gat));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n775), .B2(new_n440), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n693), .A2(G106gat), .A3(new_n426), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n769), .A2(new_n770), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT53), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n759), .A2(new_n761), .ZN(new_n785));
  INV_X1    g584(.A(new_n781), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n780), .B2(new_n787), .ZN(G1339gat));
  NOR3_X1   g587(.A1(new_n602), .A2(new_n540), .A3(new_n639), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n612), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n612), .B1(new_n631), .B2(new_n632), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n626), .A2(KEYINPUT101), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n637), .B1(new_n635), .B2(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n626), .B2(new_n612), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n627), .B2(new_n633), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n626), .A2(new_n612), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n616), .B1(new_n801), .B2(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n521), .B1(new_n519), .B2(new_n522), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n527), .A2(new_n529), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n535), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n539), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n797), .A2(new_n803), .A3(new_n634), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n571), .B1(new_n808), .B2(new_n756), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n756), .B1(new_n639), .B2(new_n807), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n797), .A2(new_n803), .A3(new_n540), .A4(new_n634), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n789), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  NOR4_X1   g612(.A1(new_n813), .A2(new_n430), .A3(new_n483), .A4(new_n486), .ZN(new_n814));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n540), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n812), .ZN(new_n816));
  INV_X1    g615(.A(new_n789), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n478), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n671), .A2(new_n649), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n204), .A3(new_n541), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n815), .A2(new_n823), .ZN(G1340gat));
  AOI21_X1  g623(.A(G120gat), .B1(new_n814), .B2(new_n639), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n822), .A2(new_n202), .A3(new_n693), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(G1341gat));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n814), .A2(new_n828), .A3(new_n571), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n212), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n814), .B2(new_n571), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n571), .A2(G127gat), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n830), .A2(new_n831), .B1(new_n822), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT117), .ZN(G1342gat));
  NAND3_X1  g633(.A1(new_n814), .A2(new_n213), .A3(new_n756), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT56), .Z(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n822), .B2(new_n601), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n818), .A2(new_n840), .A3(new_n440), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n813), .B2(new_n426), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n661), .A4(new_n821), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n541), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n661), .A2(new_n440), .A3(new_n649), .ZN(new_n845));
  AOI211_X1 g644(.A(new_n430), .B(new_n845), .C1(new_n817), .C2(new_n816), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n231), .A3(new_n540), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n232), .A3(new_n639), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n818), .A2(new_n440), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n662), .B1(new_n852), .B2(KEYINPUT57), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(new_n639), .A3(new_n821), .A4(new_n841), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n854), .B2(G148gat), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n851), .B(G148gat), .C1(new_n843), .C2(new_n693), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n850), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT119), .B(new_n850), .C1(new_n855), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1345gat));
  OAI21_X1  g661(.A(G155gat), .B1(new_n843), .B2(new_n694), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n236), .A3(new_n571), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1346gat));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n237), .A3(new_n756), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT120), .B1(new_n843), .B2(new_n601), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G162gat), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n843), .A2(KEYINPUT120), .A3(new_n601), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n671), .A2(new_n649), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n813), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n819), .ZN(new_n874));
  INV_X1    g673(.A(G169gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n874), .A2(new_n875), .A3(new_n541), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n813), .A2(new_n483), .A3(new_n872), .ZN(new_n877));
  AOI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n540), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(G1348gat));
  OAI21_X1  g678(.A(G176gat), .B1(new_n874), .B2(new_n693), .ZN(new_n880));
  INV_X1    g679(.A(G176gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n881), .A3(new_n639), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1349gat));
  OAI21_X1  g682(.A(G183gat), .B1(new_n874), .B2(new_n694), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n571), .A2(new_n342), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n877), .A2(KEYINPUT121), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n877), .B2(new_n885), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n884), .B(KEYINPUT123), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT60), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n884), .B(KEYINPUT122), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT60), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n819), .A3(new_n756), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G190gat), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT124), .B1(new_n895), .B2(G190gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n900), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n877), .A2(new_n343), .A3(new_n756), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n901), .B2(new_n906), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1351gat));
  NAND3_X1  g709(.A1(new_n853), .A2(new_n841), .A3(new_n871), .ZN(new_n911));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(new_n541), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n873), .A2(new_n440), .A3(new_n661), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT126), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n540), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n916), .B2(new_n912), .ZN(G1352gat));
  XNOR2_X1  g716(.A(KEYINPUT127), .B(G204gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n914), .A2(new_n693), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT62), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n911), .B2(new_n693), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1353gat));
  NAND3_X1  g721(.A1(new_n915), .A2(new_n302), .A3(new_n571), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n911), .A2(new_n694), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n924), .B2(G211gat), .ZN(new_n925));
  OAI211_X1 g724(.A(KEYINPUT63), .B(G211gat), .C1(new_n911), .C2(new_n694), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n925), .B2(new_n927), .ZN(G1354gat));
  NAND3_X1  g727(.A1(new_n915), .A2(new_n303), .A3(new_n756), .ZN(new_n929));
  OAI21_X1  g728(.A(G218gat), .B1(new_n911), .B2(new_n601), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


