

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XOR2_X1 U321 ( .A(n312), .B(n311), .Z(n541) );
  XOR2_X1 U322 ( .A(KEYINPUT6), .B(G148GAT), .Z(n290) );
  XNOR2_X1 U323 ( .A(G127GAT), .B(G57GAT), .ZN(n289) );
  XNOR2_X1 U324 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U325 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n292) );
  XNOR2_X1 U326 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n291) );
  XNOR2_X1 U327 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U328 ( .A(n294), .B(n293), .Z(n306) );
  XOR2_X1 U329 ( .A(G155GAT), .B(KEYINPUT3), .Z(n296) );
  XNOR2_X1 U330 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n295) );
  XNOR2_X1 U331 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U332 ( .A(KEYINPUT92), .B(n297), .Z(n397) );
  INV_X1 U333 ( .A(n397), .ZN(n304) );
  XOR2_X1 U334 ( .A(G85GAT), .B(G162GAT), .Z(n299) );
  XNOR2_X1 U335 ( .A(G29GAT), .B(G1GAT), .ZN(n298) );
  XNOR2_X1 U336 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U337 ( .A(KEYINPUT94), .B(n300), .Z(n302) );
  NAND2_X1 U338 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U339 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U340 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U341 ( .A(n306), .B(n305), .ZN(n312) );
  XNOR2_X1 U342 ( .A(KEYINPUT82), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U343 ( .A(n307), .B(G120GAT), .ZN(n308) );
  XOR2_X1 U344 ( .A(n308), .B(KEYINPUT83), .Z(n310) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XOR2_X1 U346 ( .A(n310), .B(n309), .Z(n412) );
  INV_X1 U347 ( .A(n412), .ZN(n311) );
  XOR2_X1 U348 ( .A(G113GAT), .B(G15GAT), .Z(n314) );
  XNOR2_X1 U349 ( .A(G50GAT), .B(G36GAT), .ZN(n313) );
  XNOR2_X1 U350 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U351 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n316) );
  XNOR2_X1 U352 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n315) );
  XNOR2_X1 U353 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U354 ( .A(n318), .B(n317), .ZN(n328) );
  XNOR2_X1 U355 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n319) );
  XNOR2_X1 U356 ( .A(n319), .B(G22GAT), .ZN(n376) );
  XOR2_X1 U357 ( .A(G169GAT), .B(G8GAT), .Z(n426) );
  XOR2_X1 U358 ( .A(n376), .B(n426), .Z(n321) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U360 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U361 ( .A(n322), .B(G141GAT), .Z(n326) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G43GAT), .Z(n324) );
  XNOR2_X1 U363 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n323) );
  XNOR2_X1 U364 ( .A(n324), .B(n323), .ZN(n359) );
  XNOR2_X1 U365 ( .A(n359), .B(G197GAT), .ZN(n325) );
  XNOR2_X1 U366 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U367 ( .A(n328), .B(n327), .Z(n565) );
  INV_X1 U368 ( .A(n565), .ZN(n506) );
  XOR2_X1 U369 ( .A(KEYINPUT33), .B(KEYINPUT77), .Z(n330) );
  XNOR2_X1 U370 ( .A(KEYINPUT31), .B(KEYINPUT71), .ZN(n329) );
  XNOR2_X1 U371 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U372 ( .A(n331), .B(G204GAT), .Z(n333) );
  XOR2_X1 U373 ( .A(G176GAT), .B(G64GAT), .Z(n425) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(n425), .ZN(n332) );
  XNOR2_X1 U375 ( .A(n333), .B(n332), .ZN(n344) );
  XOR2_X1 U376 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n335) );
  NAND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U378 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U379 ( .A(n336), .B(KEYINPUT75), .Z(n342) );
  XOR2_X1 U380 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n338) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n337) );
  XNOR2_X1 U382 ( .A(n338), .B(n337), .ZN(n375) );
  XOR2_X1 U383 ( .A(KEYINPUT72), .B(G78GAT), .Z(n340) );
  XNOR2_X1 U384 ( .A(G148GAT), .B(G106GAT), .ZN(n339) );
  XNOR2_X1 U385 ( .A(n340), .B(n339), .ZN(n382) );
  XNOR2_X1 U386 ( .A(n375), .B(n382), .ZN(n341) );
  XNOR2_X1 U387 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U388 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U389 ( .A(KEYINPUT73), .B(G92GAT), .Z(n346) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(KEYINPUT74), .ZN(n345) );
  XNOR2_X1 U391 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U392 ( .A(G85GAT), .B(n347), .ZN(n358) );
  XNOR2_X1 U393 ( .A(n348), .B(n358), .ZN(n570) );
  NOR2_X1 U394 ( .A1(n506), .A2(n570), .ZN(n459) );
  XOR2_X1 U395 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n350) );
  XNOR2_X1 U396 ( .A(KEYINPUT64), .B(KEYINPUT11), .ZN(n349) );
  XNOR2_X1 U397 ( .A(n350), .B(n349), .ZN(n363) );
  XOR2_X1 U398 ( .A(G50GAT), .B(G162GAT), .Z(n383) );
  XOR2_X1 U399 ( .A(G106GAT), .B(KEYINPUT10), .Z(n352) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U402 ( .A(n383), .B(n353), .Z(n355) );
  NAND2_X1 U403 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n355), .B(n354), .ZN(n357) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G190GAT), .ZN(n356) );
  XNOR2_X1 U406 ( .A(n356), .B(KEYINPUT78), .ZN(n420) );
  XOR2_X1 U407 ( .A(n357), .B(n420), .Z(n361) );
  XOR2_X1 U408 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U409 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U410 ( .A(n363), .B(n362), .ZN(n556) );
  INV_X1 U411 ( .A(n556), .ZN(n500) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G127GAT), .Z(n408) );
  XOR2_X1 U413 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n365) );
  XNOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U416 ( .A(n408), .B(n366), .Z(n368) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n368), .B(n367), .ZN(n380) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(G155GAT), .Z(n370) );
  XNOR2_X1 U420 ( .A(G8GAT), .B(G183GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U422 ( .A(G211GAT), .B(KEYINPUT14), .Z(n372) );
  XNOR2_X1 U423 ( .A(G78GAT), .B(KEYINPUT15), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U425 ( .A(n374), .B(n373), .Z(n378) );
  XNOR2_X1 U426 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U427 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U428 ( .A(n380), .B(n379), .Z(n573) );
  NAND2_X1 U429 ( .A1(n500), .A2(n573), .ZN(n381) );
  XOR2_X1 U430 ( .A(KEYINPUT16), .B(n381), .Z(n445) );
  XOR2_X1 U431 ( .A(KEYINPUT24), .B(n382), .Z(n385) );
  XNOR2_X1 U432 ( .A(G22GAT), .B(n383), .ZN(n384) );
  XNOR2_X1 U433 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U434 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n387) );
  NAND2_X1 U435 ( .A1(G228GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U436 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U437 ( .A(n389), .B(n388), .Z(n396) );
  XOR2_X1 U438 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n391) );
  XNOR2_X1 U439 ( .A(G218GAT), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U440 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U441 ( .A(n392), .B(KEYINPUT90), .Z(n394) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(G204GAT), .ZN(n393) );
  XNOR2_X1 U443 ( .A(n394), .B(n393), .ZN(n423) );
  XNOR2_X1 U444 ( .A(n423), .B(KEYINPUT93), .ZN(n395) );
  XNOR2_X1 U445 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U446 ( .A(n398), .B(n397), .Z(n543) );
  XOR2_X1 U447 ( .A(n543), .B(KEYINPUT28), .Z(n495) );
  INV_X1 U448 ( .A(n495), .ZN(n516) );
  XOR2_X1 U449 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n400) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(G176GAT), .ZN(n399) );
  XNOR2_X1 U451 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U452 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n402) );
  XNOR2_X1 U453 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U455 ( .A(n404), .B(n403), .Z(n414) );
  XOR2_X1 U456 ( .A(G71GAT), .B(G190GAT), .Z(n406) );
  XNOR2_X1 U457 ( .A(G43GAT), .B(G99GAT), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U459 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U460 ( .A1(G227GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U462 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U463 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U464 ( .A(KEYINPUT19), .B(G183GAT), .Z(n416) );
  XNOR2_X1 U465 ( .A(KEYINPUT86), .B(KEYINPUT17), .ZN(n415) );
  XNOR2_X1 U466 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U467 ( .A(KEYINPUT18), .B(n417), .Z(n419) );
  XOR2_X2 U468 ( .A(n418), .B(n419), .Z(n546) );
  INV_X1 U469 ( .A(n419), .ZN(n430) );
  XOR2_X1 U470 ( .A(n420), .B(G92GAT), .Z(n422) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U472 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U473 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U474 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U475 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U476 ( .A(n430), .B(n429), .Z(n539) );
  XOR2_X1 U477 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n431) );
  XNOR2_X1 U478 ( .A(n539), .B(n431), .ZN(n513) );
  NAND2_X1 U479 ( .A1(n546), .A2(n513), .ZN(n432) );
  NOR2_X1 U480 ( .A1(n516), .A2(n432), .ZN(n433) );
  NOR2_X1 U481 ( .A1(n541), .A2(n433), .ZN(n444) );
  XOR2_X1 U482 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n435) );
  NAND2_X1 U483 ( .A1(n543), .A2(n546), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U485 ( .A(KEYINPUT97), .B(n436), .Z(n528) );
  NAND2_X1 U486 ( .A1(n513), .A2(n528), .ZN(n437) );
  NAND2_X1 U487 ( .A1(n541), .A2(n437), .ZN(n442) );
  NOR2_X1 U488 ( .A1(n546), .A2(n539), .ZN(n438) );
  NOR2_X1 U489 ( .A1(n543), .A2(n438), .ZN(n439) );
  XNOR2_X1 U490 ( .A(KEYINPUT25), .B(n439), .ZN(n440) );
  XNOR2_X1 U491 ( .A(KEYINPUT99), .B(n440), .ZN(n441) );
  NOR2_X1 U492 ( .A1(n442), .A2(n441), .ZN(n443) );
  NOR2_X1 U493 ( .A1(n444), .A2(n443), .ZN(n454) );
  NAND2_X1 U494 ( .A1(n445), .A2(n454), .ZN(n446) );
  XOR2_X1 U495 ( .A(n446), .B(KEYINPUT100), .Z(n470) );
  NAND2_X1 U496 ( .A1(n459), .A2(n470), .ZN(n452) );
  NOR2_X1 U497 ( .A1(n541), .A2(n452), .ZN(n447) );
  XOR2_X1 U498 ( .A(n447), .B(KEYINPUT34), .Z(n448) );
  XNOR2_X1 U499 ( .A(G1GAT), .B(n448), .ZN(G1324GAT) );
  NOR2_X1 U500 ( .A1(n539), .A2(n452), .ZN(n449) );
  XOR2_X1 U501 ( .A(G8GAT), .B(n449), .Z(G1325GAT) );
  NOR2_X1 U502 ( .A1(n546), .A2(n452), .ZN(n451) );
  XNOR2_X1 U503 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(G1326GAT) );
  NOR2_X1 U505 ( .A1(n495), .A2(n452), .ZN(n453) );
  XOR2_X1 U506 ( .A(G22GAT), .B(n453), .Z(G1327GAT) );
  XNOR2_X1 U507 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n462) );
  XOR2_X1 U508 ( .A(KEYINPUT36), .B(n500), .Z(n575) );
  NAND2_X1 U509 ( .A1(n575), .A2(n454), .ZN(n455) );
  NOR2_X1 U510 ( .A1(n573), .A2(n455), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n456) );
  XOR2_X1 U512 ( .A(n457), .B(n456), .Z(n485) );
  INV_X1 U513 ( .A(n485), .ZN(n458) );
  NAND2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT38), .ZN(n468) );
  NOR2_X1 U516 ( .A1(n541), .A2(n468), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n462), .B(n461), .ZN(G1328GAT) );
  NOR2_X1 U518 ( .A1(n468), .A2(n539), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT102), .B(n463), .Z(n464) );
  XNOR2_X1 U520 ( .A(G36GAT), .B(n464), .ZN(G1329GAT) );
  XNOR2_X1 U521 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n546), .A2(n468), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(G43GAT), .B(n467), .ZN(G1330GAT) );
  NOR2_X1 U525 ( .A1(n495), .A2(n468), .ZN(n469) );
  XOR2_X1 U526 ( .A(G50GAT), .B(n469), .Z(G1331GAT) );
  INV_X1 U527 ( .A(n470), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT41), .B(n570), .Z(n548) );
  NAND2_X1 U529 ( .A1(n506), .A2(n548), .ZN(n484) );
  NOR2_X1 U530 ( .A1(n471), .A2(n484), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT105), .B(n472), .ZN(n480) );
  NOR2_X1 U532 ( .A1(n541), .A2(n480), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U535 ( .A(G57GAT), .B(n475), .Z(G1332GAT) );
  NOR2_X1 U536 ( .A1(n539), .A2(n480), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT106), .B(n476), .Z(n477) );
  XNOR2_X1 U538 ( .A(G64GAT), .B(n477), .ZN(G1333GAT) );
  NOR2_X1 U539 ( .A1(n546), .A2(n480), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(G1334GAT) );
  NOR2_X1 U542 ( .A1(n495), .A2(n480), .ZN(n482) );
  XNOR2_X1 U543 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G78GAT), .B(n483), .ZN(G1335GAT) );
  NOR2_X1 U546 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT109), .B(n486), .ZN(n494) );
  NOR2_X1 U548 ( .A1(n541), .A2(n494), .ZN(n487) );
  XOR2_X1 U549 ( .A(G85GAT), .B(n487), .Z(G1336GAT) );
  NOR2_X1 U550 ( .A1(n539), .A2(n494), .ZN(n488) );
  XOR2_X1 U551 ( .A(KEYINPUT110), .B(n488), .Z(n489) );
  XNOR2_X1 U552 ( .A(G92GAT), .B(n489), .ZN(G1337GAT) );
  NOR2_X1 U553 ( .A1(n546), .A2(n494), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1338GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n493) );
  XNOR2_X1 U557 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n493), .B(n492), .ZN(n497) );
  NOR2_X1 U559 ( .A1(n495), .A2(n494), .ZN(n496) );
  XOR2_X1 U560 ( .A(n497), .B(n496), .Z(G1339GAT) );
  AND2_X1 U561 ( .A1(n565), .A2(n548), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT46), .ZN(n499) );
  NOR2_X1 U563 ( .A1(n573), .A2(n499), .ZN(n501) );
  NAND2_X1 U564 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT47), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT114), .B(n503), .ZN(n510) );
  XOR2_X1 U567 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n505) );
  NAND2_X1 U568 ( .A1(n573), .A2(n575), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n507), .A2(n506), .ZN(n508) );
  NOR2_X1 U571 ( .A1(n570), .A2(n508), .ZN(n509) );
  NOR2_X1 U572 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT48), .ZN(n538) );
  NOR2_X1 U574 ( .A1(n541), .A2(n538), .ZN(n512) );
  NAND2_X1 U575 ( .A1(n513), .A2(n512), .ZN(n529) );
  NOR2_X1 U576 ( .A1(n546), .A2(n529), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT115), .ZN(n515) );
  NOR2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n524), .A2(n565), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G113GAT), .B(n517), .ZN(G1340GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n519) );
  NAND2_X1 U582 ( .A1(n524), .A2(n548), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n521) );
  XOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT117), .Z(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1341GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n573), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT50), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G127GAT), .B(n523), .ZN(G1342GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U590 ( .A1(n524), .A2(n556), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G134GAT), .B(n527), .ZN(G1343GAT) );
  XOR2_X1 U593 ( .A(G141GAT), .B(KEYINPUT119), .Z(n531) );
  INV_X1 U594 ( .A(n528), .ZN(n563) );
  NOR2_X1 U595 ( .A1(n529), .A2(n563), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n536), .A2(n565), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1344GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n533) );
  NAND2_X1 U599 ( .A1(n536), .A2(n548), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(n534), .ZN(G1345GAT) );
  NAND2_X1 U602 ( .A1(n536), .A2(n573), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n535), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U604 ( .A1(n556), .A2(n536), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(KEYINPUT54), .B(n540), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n564) );
  NOR2_X1 U609 ( .A1(n543), .A2(n564), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(KEYINPUT55), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n565), .A2(n557), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U614 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n552) );
  XOR2_X1 U615 ( .A(G176GAT), .B(KEYINPUT56), .Z(n550) );
  NAND2_X1 U616 ( .A1(n557), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1349GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n554) );
  NAND2_X1 U620 ( .A1(n557), .A2(n573), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G183GAT), .B(n555), .ZN(G1350GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n559) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n569) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .Z(n567) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

