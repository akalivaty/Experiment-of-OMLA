//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  XNOR2_X1  g001(.A(G104), .B(G107), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n189), .A4(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n191), .A2(G107), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(G104), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT76), .B(G101), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n190), .A2(new_n197), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n203), .B(new_n205), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n201), .A2(new_n212), .A3(KEYINPUT10), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G101), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT0), .A4(G128), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n214), .A2(new_n222), .A3(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n190), .A2(new_n197), .A3(new_n200), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n211), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT11), .A3(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n232), .A3(new_n236), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n213), .A2(new_n224), .A3(new_n227), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n201), .A2(new_n212), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n226), .A2(new_n211), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT12), .B1(new_n243), .B2(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n245), .B(new_n239), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G110), .B(G140), .ZN(new_n248));
  INV_X1    g062(.A(G227), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G953), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n213), .A2(new_n224), .A3(new_n227), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n238), .A2(KEYINPUT77), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(KEYINPUT77), .A3(new_n238), .ZN(new_n257));
  INV_X1    g071(.A(new_n251), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n252), .A2(G469), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G469), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n243), .A2(new_n238), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n245), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n243), .A2(KEYINPUT12), .A3(new_n238), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(KEYINPUT78), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n244), .B2(new_n246), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n240), .A2(new_n258), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n240), .A2(KEYINPUT79), .A3(new_n258), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n271), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n256), .A2(new_n257), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n251), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n261), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G221), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT9), .B(G234), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n262), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT80), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n286));
  INV_X1    g100(.A(new_n284), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n279), .A2(new_n261), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n265), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G214), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G119), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n292), .B2(G119), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n297), .A2(KEYINPUT66), .A3(G116), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT5), .B(new_n294), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G113), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT66), .B1(new_n297), .B2(G116), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n295), .A2(new_n292), .A3(G119), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n293), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n300), .A2(KEYINPUT2), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT81), .B1(new_n312), .B2(new_n226), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n299), .A2(new_n302), .B1(new_n306), .B2(new_n310), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n201), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n305), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n294), .ZN(new_n318));
  INV_X1    g132(.A(new_n310), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n311), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n216), .A3(new_n223), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G110), .B(G122), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n313), .A2(new_n324), .A3(new_n316), .A4(new_n322), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT6), .A4(new_n328), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n317), .A2(new_n294), .A3(new_n310), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n310), .B1(new_n317), .B2(new_n294), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n223), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n315), .B1(new_n201), .B2(new_n314), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n324), .B1(new_n336), .B2(new_n316), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(KEYINPUT6), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n323), .A2(new_n340), .A3(new_n325), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT82), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n329), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n211), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n220), .A2(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n348), .A2(G224), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n343), .A2(KEYINPUT83), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(KEYINPUT7), .B2(new_n349), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n201), .B(new_n314), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n324), .B(KEYINPUT8), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n349), .A2(KEYINPUT7), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n352), .A2(new_n328), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n262), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n350), .ZN(new_n362));
  OAI211_X1 g176(.A(KEYINPUT82), .B(new_n341), .C1(new_n337), .C2(new_n338), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n329), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT83), .ZN(new_n365));
  OAI21_X1  g179(.A(G210), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n361), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n359), .B1(new_n364), .B2(KEYINPUT83), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n343), .A2(new_n350), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n366), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n291), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n290), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n221), .A2(new_n238), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT67), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n220), .B1(new_n237), .B2(new_n235), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT67), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n383));
  XNOR2_X1  g197(.A(G134), .B(G137), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n236), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n229), .A2(G137), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n231), .A2(G134), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT65), .B(G131), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n237), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT68), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT68), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n385), .A2(new_n391), .A3(new_n388), .A4(new_n237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n392), .A3(new_n212), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n376), .B1(new_n382), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT64), .ZN(new_n395));
  OAI22_X1  g209(.A1(new_n379), .A2(new_n395), .B1(new_n389), .B2(new_n211), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n221), .A2(new_n238), .A3(new_n395), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n321), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n321), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n380), .B1(new_n221), .B2(new_n238), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n221), .A2(new_n238), .A3(new_n380), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n393), .B(new_n400), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(KEYINPUT69), .A2(G237), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT69), .A2(G237), .ZN(new_n405));
  AOI21_X1  g219(.A(G953), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G210), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT27), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G101), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n399), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n403), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n377), .A2(KEYINPUT64), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n379), .A2(new_n395), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n389), .A2(new_n211), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n376), .A4(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n211), .B1(new_n389), .B2(KEYINPUT68), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n378), .A2(new_n381), .B1(new_n419), .B2(new_n392), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n420), .B2(new_n376), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n421), .B2(new_n321), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT70), .A3(new_n410), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n413), .A2(KEYINPUT31), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n410), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n414), .B(new_n425), .C1(new_n421), .C2(new_n321), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT31), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT28), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n379), .B1(new_n419), .B2(new_n392), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(KEYINPUT71), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n400), .B1(new_n429), .B2(KEYINPUT71), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n321), .B1(new_n396), .B2(new_n397), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n403), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT28), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n426), .A2(new_n427), .B1(new_n436), .B2(new_n425), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G472), .A2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n439), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n424), .B2(new_n437), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n403), .A2(KEYINPUT73), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT73), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n420), .A2(new_n447), .A3(new_n400), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n393), .B1(new_n402), .B2(new_n401), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n449), .A2(KEYINPUT74), .A3(new_n321), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT74), .B1(new_n449), .B2(new_n321), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n446), .B(new_n448), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT28), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT29), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n425), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n432), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n432), .A2(new_n435), .A3(new_n410), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n454), .C1(new_n422), .C2(new_n410), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n262), .A3(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n445), .A2(KEYINPUT32), .B1(new_n459), .B2(G472), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT72), .B1(new_n445), .B2(KEYINPUT32), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n443), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT75), .B(G217), .Z(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(G234), .B2(new_n262), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT25), .ZN(new_n466));
  XNOR2_X1  g280(.A(G125), .B(G140), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT16), .ZN(new_n468));
  INV_X1    g282(.A(G140), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G125), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n470), .A2(KEYINPUT16), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n202), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(G146), .A3(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT23), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n297), .B2(G128), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n478), .C1(G119), .C2(new_n209), .ZN(new_n479));
  XNOR2_X1  g293(.A(G119), .B(G128), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT24), .B(G110), .Z(new_n481));
  AOI22_X1  g295(.A1(new_n479), .A2(G110), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  OAI22_X1  g297(.A1(new_n479), .A2(G110), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n467), .A2(new_n202), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n474), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT22), .B(G137), .ZN(new_n488));
  INV_X1    g302(.A(G234), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n281), .A2(new_n489), .A3(G953), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n488), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n483), .A2(new_n486), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n466), .B1(new_n496), .B2(G902), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(KEYINPUT25), .A3(new_n262), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n465), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n464), .A2(G902), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT69), .B(G237), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(G214), .A3(new_n348), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n204), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n406), .A2(G143), .A3(G214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(KEYINPUT18), .A2(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n344), .A2(G140), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n470), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n467), .A2(KEYINPUT84), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(G146), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n485), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT18), .A2(G131), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n507), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n236), .B1(new_n506), .B2(new_n507), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n474), .A3(new_n473), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n506), .A2(new_n236), .A3(new_n507), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n524), .A2(new_n521), .A3(KEYINPUT17), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n191), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n528), .B(new_n520), .C1(new_n523), .C2(new_n525), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n503), .B1(new_n532), .B2(G902), .ZN(new_n533));
  INV_X1    g347(.A(G475), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n530), .B2(new_n531), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(KEYINPUT86), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT19), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(new_n202), .C1(KEYINPUT19), .C2(new_n512), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n474), .B(new_n540), .C1(new_n524), .C2(new_n521), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n520), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n529), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n531), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n542), .B2(new_n529), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n542), .A2(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT85), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n531), .A3(new_n544), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n538), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n537), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n292), .A2(G122), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G116), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n556), .A2(new_n558), .A3(new_n194), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n194), .B1(new_n556), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n204), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n209), .A2(G143), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n562), .A2(new_n563), .A3(new_n229), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n209), .B2(G143), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n563), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n562), .A2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(G134), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT87), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n565), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n556), .A2(KEYINPUT14), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n292), .A2(G122), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n556), .B1(new_n576), .B2(KEYINPUT14), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n577), .B2(KEYINPUT89), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n579), .B(new_n556), .C1(new_n576), .C2(KEYINPUT14), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n194), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n559), .A2(KEYINPUT88), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n229), .B1(new_n562), .B2(new_n563), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n582), .B1(new_n564), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n559), .A2(KEYINPUT88), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n463), .A2(G953), .A3(new_n282), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OR3_X1    g402(.A1(new_n574), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n574), .B2(new_n586), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT90), .B(new_n588), .C1(new_n574), .C2(new_n586), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n262), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n592), .A2(new_n262), .A3(new_n593), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n555), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G952), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G953), .ZN(new_n603));
  INV_X1    g417(.A(G237), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n603), .B1(new_n489), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT21), .B(G898), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT91), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n262), .B(new_n348), .C1(G234), .C2(G237), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n601), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n375), .A2(new_n462), .A3(new_n502), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  AOI21_X1  g430(.A(G902), .B1(new_n424), .B2(new_n437), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n440), .ZN(new_n620));
  INV_X1    g434(.A(new_n502), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n285), .B2(new_n289), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT92), .Z(new_n624));
  AND2_X1   g438(.A1(new_n537), .A2(new_n554), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n592), .A2(new_n626), .A3(new_n593), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n589), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n595), .A2(G902), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n629), .A2(new_n630), .B1(new_n595), .B2(new_n594), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n612), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT93), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n374), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n367), .B1(new_n361), .B2(new_n365), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n369), .A2(new_n372), .A3(new_n366), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(KEYINPUT93), .A3(new_n291), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n633), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n554), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n548), .A2(KEYINPUT94), .A3(new_n553), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n536), .A2(new_n533), .B1(new_n597), .B2(new_n599), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n612), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n635), .B2(new_n639), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n624), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n487), .B(new_n656), .Z(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(G902), .A3(new_n464), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n499), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n613), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n375), .A2(new_n620), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AOI21_X1  g479(.A(new_n659), .B1(new_n285), .B2(new_n289), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT93), .B1(new_n638), .B2(new_n291), .ZN(new_n667));
  INV_X1    g481(.A(new_n291), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n634), .B(new_n668), .C1(new_n636), .C2(new_n637), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n462), .B(new_n666), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n610), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n605), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n548), .A2(KEYINPUT94), .A3(new_n553), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT94), .B1(new_n548), .B2(new_n553), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n649), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n648), .A2(KEYINPUT97), .A3(new_n649), .A4(new_n673), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT98), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n462), .A2(new_n666), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n635), .A2(new_n639), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .A4(new_n680), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XOR2_X1   g502(.A(new_n673), .B(KEYINPUT39), .Z(new_n689));
  OR2_X1    g503(.A1(new_n290), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n638), .B(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n413), .A2(new_n423), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n452), .A2(new_n425), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n262), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n445), .A2(KEYINPUT32), .B1(new_n700), .B2(G472), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n443), .A3(new_n461), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n600), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n625), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n291), .A3(new_n659), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n697), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n693), .A2(new_n694), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n204), .ZN(G45));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n710));
  INV_X1    g524(.A(new_n673), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n625), .A2(new_n631), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n710), .B1(new_n670), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n683), .A2(KEYINPUT101), .A3(new_n685), .A4(new_n712), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OR2_X1    g531(.A1(new_n279), .A2(new_n261), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n279), .A2(new_n261), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n287), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n462), .A2(new_n502), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n640), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n651), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND2_X1  g541(.A1(new_n660), .A2(new_n462), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n721), .B1(new_n667), .B2(new_n669), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n721), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n297), .ZN(G21));
  INV_X1    g548(.A(new_n705), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n635), .B2(new_n639), .ZN(new_n736));
  INV_X1    g550(.A(new_n424), .ZN(new_n737));
  INV_X1    g551(.A(new_n432), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n452), .B2(KEYINPUT28), .ZN(new_n739));
  OAI22_X1  g553(.A1(new_n739), .A2(new_n410), .B1(KEYINPUT31), .B2(new_n411), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n439), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(new_n502), .C1(new_n618), .C2(new_n617), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT103), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n619), .A2(new_n744), .A3(new_n502), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n720), .A2(new_n611), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n736), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  AND2_X1   g563(.A1(new_n619), .A2(new_n741), .ZN(new_n750));
  INV_X1    g564(.A(new_n659), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n713), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT102), .B1(new_n685), .B2(new_n721), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n730), .B(new_n720), .C1(new_n635), .C2(new_n639), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  AOI21_X1  g571(.A(KEYINPUT104), .B1(new_n247), .B2(new_n251), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n252), .A2(new_n259), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(KEYINPUT104), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n263), .B1(new_n760), .B2(G469), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n284), .B1(new_n761), .B2(new_n719), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n636), .A2(new_n291), .A3(new_n637), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n440), .A2(new_n442), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n621), .B1(new_n460), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n767), .A3(new_n712), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT42), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(new_n765), .A3(new_n462), .A4(new_n502), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n236), .ZN(G33));
  NAND4_X1  g587(.A1(new_n680), .A2(new_n462), .A3(new_n502), .A4(new_n765), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT105), .B(G134), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G36));
  INV_X1    g590(.A(new_n631), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n625), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT43), .Z(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n751), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n620), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT44), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n760), .A2(KEYINPUT106), .A3(KEYINPUT45), .ZN(new_n785));
  INV_X1    g599(.A(new_n759), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n785), .B(G469), .C1(KEYINPUT45), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT106), .B1(new_n760), .B2(KEYINPUT45), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n264), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n288), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n287), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n689), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n782), .A2(new_n783), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n764), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n784), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n287), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n462), .A2(new_n713), .A3(new_n502), .A4(new_n764), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  OR4_X1    g619(.A1(new_n621), .A2(new_n778), .A3(new_n668), .A4(new_n284), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n718), .A2(new_n719), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT49), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n806), .A2(KEYINPUT108), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n703), .A3(new_n697), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n761), .A2(new_n719), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n499), .A2(new_n658), .A3(new_n711), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n287), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n762), .A2(KEYINPUT110), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n702), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n705), .B1(new_n667), .B2(new_n669), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n714), .B2(new_n715), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n813), .A2(new_n824), .A3(new_n687), .A4(new_n756), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n731), .A2(new_n732), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n826), .A2(new_n753), .B1(new_n682), .B2(new_n686), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n813), .B1(new_n827), .B2(new_n824), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n748), .A2(new_n723), .A3(new_n726), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT109), .B1(new_n830), .B2(new_n733), .ZN(new_n831));
  INV_X1    g645(.A(new_n728), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n754), .B2(new_n755), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n722), .B1(new_n640), .B2(new_n651), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n748), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n777), .A2(new_n625), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n611), .A3(new_n601), .ZN(new_n838));
  INV_X1    g652(.A(new_n374), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n620), .A3(new_n839), .A4(new_n622), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n615), .A2(new_n774), .A3(new_n661), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n750), .A2(new_n751), .A3(new_n712), .A4(new_n762), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n537), .A2(new_n648), .A3(new_n704), .A4(new_n673), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n462), .A2(new_n843), .A3(new_n666), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n764), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n841), .A2(new_n772), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n831), .A2(new_n836), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n829), .A2(KEYINPUT111), .A3(KEYINPUT53), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n824), .A2(new_n687), .A3(new_n756), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n827), .A2(new_n813), .A3(new_n824), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n831), .A2(new_n836), .A3(new_n846), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n825), .A3(new_n828), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT111), .B1(new_n857), .B2(KEYINPUT53), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n852), .A3(new_n851), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n830), .A2(new_n733), .A3(new_n849), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n846), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n860), .A2(new_n849), .B1(new_n829), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n859), .A2(KEYINPUT113), .A3(new_n865), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n764), .A2(new_n720), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n605), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n874), .A2(new_n502), .A3(new_n703), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n625), .A3(new_n631), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT117), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n284), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n800), .A2(new_n801), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n779), .A2(new_n606), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n746), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n764), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n874), .A2(new_n779), .ZN(new_n885));
  INV_X1    g699(.A(new_n752), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n881), .A2(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n883), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n696), .A2(new_n291), .A3(new_n720), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(KEYINPUT50), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(KEYINPUT115), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT50), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n877), .B(new_n887), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n891), .B(new_n892), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT51), .A3(new_n877), .A4(new_n887), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n885), .A2(new_n767), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT48), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n875), .A2(new_n632), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n888), .A2(new_n826), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n603), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n897), .A2(new_n899), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n868), .A2(new_n869), .A3(new_n908), .A4(KEYINPUT119), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n602), .A2(new_n348), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n851), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT111), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n855), .A3(new_n848), .ZN(new_n915));
  AOI221_X4 g729(.A(new_n867), .B1(new_n863), .B2(new_n864), .C1(new_n915), .C2(KEYINPUT54), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT113), .B1(new_n859), .B2(new_n865), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT119), .B1(new_n918), .B2(new_n908), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n812), .B1(new_n911), .B2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n863), .A2(new_n262), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(G210), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(KEYINPUT120), .A3(G210), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n343), .A2(new_n350), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n364), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT55), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(KEYINPUT56), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n921), .A2(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n931), .B2(KEYINPUT56), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n348), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n930), .A2(new_n932), .A3(new_n937), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G51));
  NAND2_X1  g753(.A1(new_n276), .A2(new_n278), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n829), .A2(new_n862), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n855), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n864), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n263), .B(KEYINPUT57), .Z(new_n944));
  OAI21_X1  g758(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n787), .A2(new_n788), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n921), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n933), .B1(new_n945), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n921), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n551), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT122), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n933), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n921), .A2(new_n954), .A3(new_n551), .A4(new_n949), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT123), .ZN(G60));
  INV_X1    g771(.A(new_n629), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  NOR3_X1   g774(.A1(new_n943), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n916), .B2(new_n917), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n933), .B(new_n961), .C1(new_n963), .C2(new_n958), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT60), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n942), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT124), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n933), .B1(new_n968), .B2(new_n496), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n657), .B(KEYINPUT125), .Z(new_n970));
  OAI211_X1 g784(.A(new_n969), .B(KEYINPUT61), .C1(new_n968), .C2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n967), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n934), .B1(new_n974), .B2(new_n495), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n968), .A2(new_n970), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n977), .ZN(G66));
  AOI21_X1  g792(.A(new_n348), .B1(new_n608), .B2(G224), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n615), .A2(new_n661), .A3(new_n840), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n831), .A2(new_n836), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n981), .B2(new_n348), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n363), .B(new_n329), .C1(G898), .C2(new_n348), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G69));
  AND2_X1   g798(.A1(new_n797), .A2(new_n804), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n827), .A2(new_n716), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n794), .A2(new_n736), .A3(new_n767), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n769), .A2(new_n771), .A3(new_n774), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n539), .B1(KEYINPUT19), .B2(new_n512), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n421), .B(new_n992), .Z(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n671), .B2(new_n348), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n708), .A2(new_n986), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n837), .A2(new_n764), .A3(new_n601), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n691), .A2(new_n462), .A3(new_n502), .A4(new_n999), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1001));
  NAND4_X1  g815(.A1(new_n997), .A2(new_n998), .A3(new_n985), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n993), .B1(new_n1002), .B2(new_n348), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n249), .B2(new_n671), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n1002), .B2(new_n981), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n422), .A2(new_n425), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1008), .B1(new_n990), .B2(new_n981), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n422), .A3(new_n425), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1013), .A3(new_n934), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n422), .A2(new_n410), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n915), .B(new_n1008), .C1(new_n698), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(G57));
endmodule


