//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT65), .B(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT66), .B(KEYINPUT1), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n209), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT67), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(KEYINPUT13), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n212), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n262), .B(new_n264), .C1(G232), .C2(new_n263), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT75), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n257), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n275), .A2(G238), .A3(new_n255), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n253), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n265), .B2(new_n270), .ZN(new_n279));
  NOR4_X1   g0079(.A1(new_n279), .A2(KEYINPUT13), .A3(new_n257), .A4(new_n276), .ZN(new_n280));
  OAI21_X1  g0080(.A(G169), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n278), .ZN(new_n285));
  INV_X1    g0085(.A(new_n280), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G179), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n288));
  OAI211_X1 g0088(.A(G169), .B(new_n282), .C1(new_n278), .C2(new_n280), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n229), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G13), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT12), .B1(new_n292), .B2(new_n222), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT77), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR3_X1    g0095(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n294), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n259), .A2(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G77), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n300), .B1(new_n211), .B2(new_n302), .C1(new_n222), .C2(new_n229), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n304), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT68), .B1(new_n304), .B2(new_n228), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(new_n228), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n254), .A2(G20), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G68), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n303), .A2(new_n307), .A3(new_n309), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n298), .A2(new_n311), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n290), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G238), .A2(G1698), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n262), .B(new_n319), .C1(new_n237), .C2(G1698), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT70), .B(G107), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n320), .B(new_n272), .C1(new_n262), .C2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n257), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n275), .A2(new_n255), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G244), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(KEYINPUT8), .A2(G58), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT8), .A2(G58), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT15), .B(G87), .Z(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n301), .B1(new_n335), .B2(new_n299), .ZN(new_n336));
  INV_X1    g0136(.A(G77), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n229), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G13), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n314), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n338), .A2(new_n312), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n313), .A2(G77), .A3(new_n314), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n330), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n327), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n299), .A2(new_n331), .A3(new_n332), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n301), .A2(G150), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n307), .B1(new_n211), .B2(new_n340), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n291), .A2(new_n211), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n292), .B(new_n352), .C1(new_n305), .C2(new_n306), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n263), .A2(G222), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G223), .A2(G1698), .ZN(new_n356));
  AND2_X1   g0156(.A1(KEYINPUT3), .A2(G33), .ZN(new_n357));
  NOR2_X1   g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n260), .A2(new_n337), .A3(new_n261), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n272), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n275), .A2(G226), .A3(new_n255), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n324), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n363), .A2(G179), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT69), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n367), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n354), .B(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n346), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n285), .A2(new_n286), .A3(G190), .ZN(new_n372));
  INV_X1    g0172(.A(new_n317), .ZN(new_n373));
  OAI21_X1  g0173(.A(G200), .B1(new_n278), .B2(new_n280), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n328), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n327), .A2(new_n364), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n343), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n318), .A2(new_n371), .A3(new_n375), .A4(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n275), .A2(G232), .A3(new_n255), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n259), .A2(new_n219), .ZN(new_n383));
  INV_X1    g0183(.A(G223), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n260), .A2(new_n261), .B1(new_n384), .B2(new_n263), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n212), .A2(G1698), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n382), .B(new_n324), .C1(new_n387), .C2(new_n275), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(G179), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(KEYINPUT80), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n263), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n386), .C1(new_n357), .C2(new_n358), .ZN(new_n392));
  INV_X1    g0192(.A(new_n383), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n257), .B1(new_n394), .B2(new_n272), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT80), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n382), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n398), .B2(new_n364), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT81), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n222), .B2(G58), .ZN(new_n405));
  INV_X1    g0205(.A(G159), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n405), .A2(new_n229), .B1(new_n406), .B2(new_n302), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n260), .A2(new_n229), .A3(new_n261), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n261), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n223), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n403), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n357), .A2(new_n358), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n414), .B2(new_n229), .ZN(new_n415));
  INV_X1    g0215(.A(new_n411), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n302), .A2(new_n406), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT65), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G68), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n421), .A3(G58), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n203), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n423), .B2(G20), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n417), .A2(new_n424), .A3(KEYINPUT16), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n413), .A2(new_n312), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n307), .A2(new_n340), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n333), .A2(new_n291), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n428), .A2(new_n429), .B1(new_n340), .B2(new_n333), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n426), .B2(new_n430), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n399), .B(new_n402), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n400), .A2(new_n401), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n388), .A2(G190), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n398), .B2(new_n329), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n425), .A2(new_n312), .ZN(new_n439));
  INV_X1    g0239(.A(new_n412), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT16), .B1(new_n440), .B2(new_n424), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n430), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n426), .A2(new_n430), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n396), .B1(new_n395), .B2(new_n382), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n275), .B1(new_n392), .B2(new_n393), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n446), .A2(KEYINPUT80), .A3(new_n381), .A4(new_n257), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n329), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n436), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT17), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n442), .A2(KEYINPUT79), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n434), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n399), .A3(new_n402), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n350), .A2(new_n307), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT9), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT71), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n340), .A2(new_n211), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n353), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n459), .A2(KEYINPUT71), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT72), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n363), .A2(G200), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n345), .B2(new_n363), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(new_n463), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT72), .ZN(new_n471));
  INV_X1    g0271(.A(new_n463), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n351), .A2(new_n460), .A3(new_n353), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT73), .B(KEYINPUT10), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n466), .A2(new_n469), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n469), .B1(new_n464), .B2(new_n465), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT74), .A3(KEYINPUT10), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT74), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n468), .B1(new_n470), .B2(new_n473), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT10), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n476), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n435), .A2(new_n452), .A3(new_n457), .A4(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n380), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n220), .A2(new_n263), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n262), .B(new_n486), .C1(G257), .C2(new_n263), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n275), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n254), .A2(G45), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  AOI211_X1 g0292(.A(new_n216), .B(new_n272), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n490), .A2(new_n256), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n364), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n496), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n489), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(G179), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n229), .A2(KEYINPUT23), .A3(G107), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT70), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n215), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT70), .A2(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n229), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n229), .B(G87), .C1(new_n357), .C2(new_n358), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT22), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n262), .A2(new_n512), .A3(new_n229), .A4(G87), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n299), .A2(G116), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n501), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n513), .ZN(new_n517));
  INV_X1    g0317(.A(new_n506), .ZN(new_n518));
  NOR2_X1   g0318(.A1(KEYINPUT70), .A2(G107), .ZN(new_n519));
  OAI21_X1  g0319(.A(G20), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n502), .B1(new_n520), .B2(KEYINPUT23), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n517), .A2(new_n501), .A3(new_n521), .A4(new_n515), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n312), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n340), .A2(new_n215), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n525), .B(KEYINPUT25), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n254), .A2(G33), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n292), .B(new_n527), .C1(new_n305), .C2(new_n306), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n215), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n524), .A2(KEYINPUT87), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT87), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n517), .A2(new_n515), .A3(new_n521), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT24), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n313), .B1(new_n534), .B2(new_n522), .ZN(new_n535));
  INV_X1    g0335(.A(new_n530), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n500), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n524), .A2(new_n530), .ZN(new_n539));
  NOR4_X1   g0339(.A1(new_n489), .A2(new_n493), .A3(new_n345), .A4(new_n498), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n499), .A2(new_n329), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(G244), .C1(new_n358), .C2(new_n357), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  INV_X1    g0347(.A(G244), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n260), .B2(new_n261), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n547), .C1(new_n549), .C2(KEYINPUT4), .ZN(new_n550));
  OAI21_X1  g0350(.A(G250), .B1(new_n357), .B2(new_n358), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n263), .B1(new_n551), .B2(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n272), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n228), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n492), .A2(new_n491), .B1(new_n554), .B2(new_n274), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(G257), .ZN(new_n557));
  AND2_X1   g0357(.A1(KEYINPUT5), .A2(G41), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT5), .A2(G41), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(new_n275), .C1(new_n560), .C2(new_n490), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n553), .A2(new_n563), .A3(new_n496), .ZN(new_n564));
  AND2_X1   g0364(.A1(KEYINPUT83), .A2(G200), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  INV_X1    g0367(.A(G97), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n215), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n229), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n322), .B1(new_n415), .B2(new_n416), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n302), .A2(new_n337), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n312), .B1(new_n568), .B2(new_n340), .ZN(new_n579));
  INV_X1    g0379(.A(new_n528), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G97), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n345), .B1(new_n329), .B2(KEYINPUT83), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n553), .A2(new_n563), .A3(new_n496), .A4(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n566), .A2(new_n579), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n564), .A2(new_n364), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n340), .A2(new_n568), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n321), .B1(new_n410), .B2(new_n411), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n587), .A2(new_n573), .A3(new_n576), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n581), .C1(new_n588), .C2(new_n313), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n553), .A2(new_n563), .A3(new_n376), .A4(new_n496), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(G238), .B(new_n263), .C1(new_n357), .C2(new_n358), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT84), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n262), .A2(new_n595), .A3(G238), .A4(new_n263), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(G33), .A2(G116), .ZN(new_n598));
  OAI211_X1 g0398(.A(G244), .B(G1698), .C1(new_n357), .C2(new_n358), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n272), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n272), .A2(new_n491), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n495), .B1(new_n602), .B2(G250), .ZN(new_n603));
  AOI21_X1  g0403(.A(G169), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n599), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n594), .B2(new_n596), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n275), .B1(new_n607), .B2(new_n598), .ZN(new_n608));
  INV_X1    g0408(.A(new_n603), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n608), .A2(G179), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n335), .A2(new_n292), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G87), .A2(G97), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n321), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT19), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n268), .B2(new_n269), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(G20), .ZN(new_n617));
  INV_X1    g0417(.A(new_n299), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n615), .B1(new_n618), .B2(new_n568), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n229), .B(G68), .C1(new_n357), .C2(new_n358), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n262), .A2(KEYINPUT85), .A3(new_n229), .A4(G68), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n617), .A2(new_n619), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n612), .B1(new_n624), .B2(new_n312), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n580), .A2(new_n335), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n605), .B(new_n611), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n263), .A2(G257), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n262), .B(new_n631), .C1(new_n216), .C2(new_n263), .ZN(new_n632));
  INV_X1    g0432(.A(G303), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n414), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n272), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n555), .A2(G270), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n496), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n376), .ZN(new_n638));
  INV_X1    g0438(.A(G116), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n340), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n313), .A2(new_n292), .A3(G116), .A4(new_n527), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n304), .A2(new_n228), .B1(G20), .B2(new_n639), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n547), .B(new_n229), .C1(G33), .C2(new_n568), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n642), .A2(KEYINPUT20), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT20), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n640), .B(new_n641), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n637), .A2(G169), .A3(new_n646), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n637), .A2(G200), .ZN(new_n651));
  INV_X1    g0451(.A(new_n646), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n635), .A2(G190), .A3(new_n496), .A4(new_n636), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n637), .A2(KEYINPUT21), .A3(G169), .A4(new_n646), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n647), .A2(new_n650), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n608), .A2(new_n609), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G190), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n624), .A2(new_n312), .ZN(new_n659));
  INV_X1    g0459(.A(new_n612), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n580), .A2(G87), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(G200), .B1(new_n608), .B2(new_n609), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n658), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n630), .A2(new_n656), .A3(new_n665), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n485), .A2(new_n543), .A3(new_n592), .A4(new_n666), .ZN(G372));
  OR4_X1    g0467(.A1(new_n535), .A2(new_n541), .A3(new_n536), .A4(new_n540), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n329), .B1(new_n601), .B2(new_n603), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n662), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n664), .A2(KEYINPUT88), .A3(new_n625), .A4(new_n661), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n658), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n668), .A2(new_n592), .A3(new_n630), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n650), .A2(new_n647), .A3(new_n655), .ZN(new_n675));
  INV_X1    g0475(.A(new_n500), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n539), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n630), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n591), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n673), .A2(new_n679), .A3(new_n630), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n630), .A2(KEYINPUT26), .A3(new_n665), .A4(new_n679), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n659), .A2(new_n660), .A3(new_n627), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT86), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n604), .A2(new_n610), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n670), .A2(new_n662), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n658), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n679), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n682), .A2(new_n685), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n485), .B1(new_n678), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n370), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n399), .A2(new_n442), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n401), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n379), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n290), .A2(new_n317), .B1(new_n375), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n452), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT90), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n483), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n476), .A2(new_n478), .A3(new_n482), .A4(KEYINPUT90), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n696), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n695), .A2(new_n709), .ZN(G369));
  NOR2_X1   g0510(.A1(new_n339), .A2(G20), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n254), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G213), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G343), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n676), .A2(new_n539), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT87), .B1(new_n524), .B2(new_n530), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n535), .A2(new_n532), .A3(new_n536), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n676), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n668), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT91), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n724), .A2(new_n726), .A3(new_n718), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT91), .B1(new_n538), .B2(new_n717), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n675), .A2(new_n718), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n720), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n717), .A2(new_n646), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n656), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n675), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n735), .B2(new_n733), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n739), .ZN(G399));
  INV_X1    g0540(.A(new_n207), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G41), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n321), .A2(new_n639), .A3(new_n613), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n742), .A2(new_n743), .A3(new_n254), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT92), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT92), .ZN(new_n746));
  INV_X1    g0546(.A(new_n742), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n745), .B(new_n746), .C1(new_n233), .C2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  AND4_X1   g0549(.A1(new_n668), .A2(new_n592), .A3(new_n630), .A4(new_n673), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT95), .B1(new_n724), .B2(new_n735), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT95), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n538), .A2(new_n752), .A3(new_n675), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n630), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n692), .A2(new_n681), .A3(new_n679), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n750), .B(KEYINPUT96), .C1(new_n751), .C2(new_n753), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n756), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(KEYINPUT29), .A3(new_n718), .ZN(new_n763));
  INV_X1    g0563(.A(new_n677), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n757), .B1(new_n750), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n682), .A2(new_n685), .A3(new_n693), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n717), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT94), .B1(new_n767), .B2(KEYINPUT29), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n718), .B1(new_n694), .B2(new_n678), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT94), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT29), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n763), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n601), .A2(new_n494), .A3(new_n603), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n638), .ZN(new_n778));
  INV_X1    g0578(.A(new_n564), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n775), .B2(new_n776), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n774), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n638), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n775), .B2(new_n776), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n657), .A2(KEYINPUT93), .A3(new_n494), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n783), .A2(KEYINPUT30), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n564), .A2(new_n376), .A3(new_n637), .ZN(new_n786));
  OR3_X1    g0586(.A1(new_n786), .A2(new_n499), .A3(new_n657), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n781), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n717), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT31), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n543), .A2(new_n666), .A3(new_n592), .A4(new_n718), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(KEYINPUT31), .A3(new_n717), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G330), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n773), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n749), .B1(new_n796), .B2(new_n254), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT97), .ZN(G364));
  AOI21_X1  g0598(.A(new_n254), .B1(new_n711), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n742), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n738), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n736), .ZN(new_n803));
  INV_X1    g0603(.A(new_n801), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n229), .A2(new_n376), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n345), .A3(new_n329), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR4_X1   g0607(.A1(new_n229), .A2(new_n376), .A3(new_n345), .A4(G200), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(G77), .B1(new_n808), .B2(G58), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT99), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n229), .A2(G190), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G179), .A2(G200), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n406), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n229), .B1(new_n812), .B2(G190), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n568), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n805), .A2(G190), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n329), .A2(G179), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n811), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n818), .A2(new_n211), .B1(new_n820), .B2(new_n215), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n805), .A2(new_n345), .A3(G200), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n817), .B(new_n821), .C1(G68), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n819), .A2(G20), .A3(G190), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n262), .B1(new_n825), .B2(new_n219), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT100), .Z(new_n827));
  NAND4_X1  g0627(.A1(new_n810), .A2(new_n815), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT101), .Z(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n414), .B1(new_n825), .B2(new_n633), .ZN(new_n832));
  INV_X1    g0632(.A(new_n813), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G329), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n818), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G311), .A2(new_n807), .B1(new_n835), .B2(G326), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT33), .B(G317), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n823), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n816), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G322), .A2(new_n808), .B1(new_n839), .B2(G294), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n834), .A2(new_n836), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n829), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n228), .B1(G20), .B2(new_n364), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n804), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n233), .A2(G45), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n248), .A2(G45), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n741), .A2(new_n262), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n847), .C2(new_n846), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n741), .A2(new_n414), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G355), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(G116), .C2(new_n207), .ZN(new_n853));
  NOR2_X1   g0653(.A1(G13), .A2(G33), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(G20), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n843), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n856), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n844), .B(new_n858), .C1(new_n736), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n803), .A2(new_n860), .ZN(G396));
  NAND2_X1  g0661(.A1(new_n343), .A2(new_n717), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n346), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n379), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n701), .A2(new_n718), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n769), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n718), .B(new_n868), .C1(new_n694), .C2(new_n678), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n795), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n804), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n843), .A2(new_n854), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n801), .B1(new_n875), .B2(G77), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT102), .ZN(new_n877));
  INV_X1    g0677(.A(new_n843), .ZN(new_n878));
  INV_X1    g0678(.A(G132), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n262), .B1(new_n813), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n820), .A2(new_n202), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n201), .B2(new_n816), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n823), .A2(G150), .B1(new_n808), .B2(G143), .ZN(new_n884));
  INV_X1    g0684(.A(G137), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n884), .B1(new_n885), .B2(new_n818), .C1(new_n406), .C2(new_n806), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT34), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n888), .B1(new_n887), .B2(new_n886), .C1(new_n211), .C2(new_n825), .ZN(new_n889));
  INV_X1    g0689(.A(new_n808), .ZN(new_n890));
  INV_X1    g0690(.A(G294), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n890), .A2(new_n891), .B1(new_n830), .B2(new_n822), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(G303), .B2(new_n835), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n833), .A2(G311), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n817), .B1(G116), .B2(new_n807), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n820), .A2(new_n219), .ZN(new_n896));
  INV_X1    g0696(.A(new_n825), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n262), .B(new_n896), .C1(G107), .C2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n877), .B1(new_n878), .B2(new_n900), .C1(new_n868), .C2(new_n855), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n873), .A2(new_n901), .ZN(G384));
  NAND3_X1  g0702(.A1(new_n435), .A2(new_n452), .A3(new_n457), .ZN(new_n903));
  INV_X1    g0703(.A(new_n715), .ZN(new_n904));
  INV_X1    g0704(.A(new_n430), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT16), .B1(new_n417), .B2(new_n424), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n906), .A2(new_n306), .A3(new_n305), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n425), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n399), .A2(new_n904), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT37), .B1(new_n912), .B2(new_n455), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n444), .A2(new_n450), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n911), .B2(new_n908), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n910), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n373), .A2(new_n718), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n318), .A2(new_n375), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n375), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n317), .B(new_n717), .C1(new_n927), .C2(new_n290), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n868), .ZN(new_n930));
  NOR2_X1   g0730(.A1(KEYINPUT105), .A2(KEYINPUT31), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n788), .A2(new_n717), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n792), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n932), .B1(new_n788), .B2(new_n717), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n930), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n923), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n904), .B1(new_n431), .B2(new_n432), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n914), .A3(new_n697), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n913), .A2(new_n914), .B1(new_n943), .B2(KEYINPUT37), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n700), .B2(new_n452), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n920), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n922), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(KEYINPUT40), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT106), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n485), .B1(new_n934), .B2(new_n936), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n950), .B(new_n951), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(G330), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT39), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n921), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n318), .A2(new_n717), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n698), .A2(new_n699), .A3(new_n715), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n869), .A2(new_n865), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n923), .A3(new_n929), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT104), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT104), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n961), .A3(new_n964), .A4(new_n959), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n953), .B(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n763), .A2(new_n485), .A3(new_n768), .A4(new_n772), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n709), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n254), .B2(new_n711), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n571), .A2(new_n572), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT103), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n639), .B1(new_n973), .B2(KEYINPUT35), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n230), .C1(KEYINPUT35), .C2(new_n973), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT36), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n422), .A2(G77), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n233), .A2(new_n977), .B1(G50), .B2(new_n202), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(G1), .A3(new_n339), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n971), .A2(new_n976), .A3(new_n979), .ZN(G367));
  INV_X1    g0780(.A(new_n820), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(G97), .ZN(new_n982));
  INV_X1    g0782(.A(G317), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n414), .C1(new_n983), .C2(new_n813), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n822), .A2(new_n891), .B1(new_n816), .B2(new_n321), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT46), .B1(new_n897), .B2(G116), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n830), .B2(new_n806), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT110), .B(G311), .Z(new_n989));
  AOI22_X1  g0789(.A1(new_n835), .A2(new_n989), .B1(new_n808), .B2(G303), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT111), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n897), .A2(KEYINPUT46), .A3(G116), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT112), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n988), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n897), .A2(G58), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n807), .A2(G50), .B1(new_n808), .B2(G150), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n202), .B2(new_n816), .ZN(new_n997));
  INV_X1    g0797(.A(G143), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n998), .A2(new_n818), .B1(new_n822), .B2(new_n406), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n262), .B1(new_n813), .B2(new_n885), .C1(new_n337), .C2(new_n820), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n994), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT47), .Z(new_n1003));
  AOI21_X1  g0803(.A(new_n804), .B1(new_n1003), .B2(new_n843), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n335), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n849), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n857), .B1(new_n207), .B2(new_n1005), .C1(new_n244), .C2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n757), .A2(new_n662), .A3(new_n717), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n673), .B(new_n630), .C1(new_n663), .C2(new_n718), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1004), .B(new_n1007), .C1(new_n859), .C2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n589), .A2(new_n717), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n592), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n679), .A2(new_n717), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n739), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT43), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n591), .B1(new_n1013), .B2(new_n724), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT107), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT107), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n591), .C1(new_n1013), .C2(new_n724), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n718), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1015), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n729), .A2(new_n731), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT42), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n726), .B1(new_n724), .B2(new_n718), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n538), .A2(KEYINPUT91), .A3(new_n717), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n730), .B1(new_n1031), .B2(new_n725), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(KEYINPUT42), .A3(new_n1025), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1024), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1010), .B1(new_n1034), .B2(KEYINPUT108), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT42), .B1(new_n1032), .B2(new_n1025), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1029), .A2(new_n1030), .B1(new_n543), .B2(new_n723), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1037), .A2(new_n1027), .A3(new_n730), .A4(new_n1015), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1023), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT108), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1010), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1018), .B(new_n1034), .C1(new_n1035), .C2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1035), .A2(new_n1042), .A3(new_n1018), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1017), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(KEYINPUT43), .A3(new_n1039), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n1016), .A3(new_n1044), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n799), .B(KEYINPUT109), .Z(new_n1051));
  AND2_X1   g0851(.A1(new_n768), .A2(new_n772), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n871), .B1(new_n1052), .B2(new_n763), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n739), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n719), .B(new_n1025), .C1(new_n1037), .C2(new_n730), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT45), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT44), .B1(new_n732), .B2(new_n1025), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT44), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n1015), .C1(new_n1032), .C2(new_n720), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1054), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT45), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1055), .B(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1063), .A2(new_n739), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1037), .B(new_n730), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(new_n738), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1053), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n742), .B(KEYINPUT41), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1051), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1011), .B1(new_n1050), .B2(new_n1071), .ZN(G387));
  AOI21_X1  g0872(.A(new_n1006), .B1(new_n240), .B2(G45), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n743), .B2(new_n851), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n334), .A2(new_n211), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT50), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n202), .A2(new_n337), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1076), .A2(G45), .A3(new_n743), .A4(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1074), .A2(new_n1078), .B1(G107), .B2(new_n207), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n804), .B1(new_n1079), .B2(new_n857), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n202), .A2(new_n806), .B1(new_n822), .B2(new_n333), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT113), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n897), .A2(G77), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n833), .A2(G150), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1083), .A2(new_n982), .A3(new_n1084), .A4(new_n262), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n890), .A2(new_n211), .B1(new_n1005), .B2(new_n816), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1082), .B(new_n1087), .C1(new_n406), .C2(new_n818), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G303), .A2(new_n807), .B1(new_n835), .B2(G322), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n983), .B2(new_n890), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n823), .B2(new_n989), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n830), .B2(new_n816), .C1(new_n891), .C2(new_n825), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n262), .B1(new_n833), .B2(G326), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n820), .A2(new_n639), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1088), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT114), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1080), .B1(new_n729), .B2(new_n859), .C1(new_n1102), .C2(new_n878), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1067), .A2(new_n1051), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1068), .A2(new_n796), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1067), .A2(new_n773), .A3(new_n795), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n742), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(G393));
  OAI221_X1 g0909(.A(new_n857), .B1(new_n568), .B2(new_n207), .C1(new_n251), .C2(new_n1006), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n835), .A2(G317), .B1(new_n808), .B2(G311), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT52), .Z(new_n1112));
  OAI22_X1  g0912(.A1(new_n822), .A2(new_n633), .B1(new_n816), .B2(new_n639), .ZN(new_n1113));
  INV_X1    g0913(.A(G322), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n414), .B1(new_n813), .B2(new_n1114), .C1(new_n215), .C2(new_n820), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(G283), .C2(new_n897), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1112), .B(new_n1116), .C1(new_n891), .C2(new_n806), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n807), .A2(new_n334), .B1(new_n839), .B2(G77), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n211), .B2(new_n822), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1119), .A2(KEYINPUT115), .ZN(new_n1120));
  INV_X1    g0920(.A(G150), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n890), .A2(new_n406), .B1(new_n818), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(KEYINPUT115), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n414), .B(new_n896), .C1(G143), .C2(new_n833), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n223), .A2(new_n825), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1117), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n804), .B1(new_n1128), .B2(new_n843), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1110), .B(new_n1129), .C1(new_n1025), .C2(new_n859), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1051), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1065), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1053), .A2(new_n1064), .A3(new_n1061), .A4(new_n1067), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n747), .B1(new_n1065), .B2(new_n1107), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G390));
  AND3_X1   g0936(.A1(new_n864), .A2(G330), .A3(new_n865), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n934), .B2(new_n936), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n929), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n957), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n947), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n762), .A2(new_n718), .A3(new_n864), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n865), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n929), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1139), .B1(new_n869), .B2(new_n865), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(new_n1142), .B1(new_n955), .B2(new_n956), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1141), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n955), .A2(new_n956), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n957), .B2(new_n1147), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n794), .A2(new_n929), .A3(new_n1137), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1139), .B1(new_n1144), .B2(new_n865), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1152), .B(new_n1154), .C1(new_n1155), .C2(new_n1143), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1144), .A2(new_n865), .A3(new_n1153), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n929), .B1(new_n794), .B2(new_n1137), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n960), .B1(new_n1140), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n485), .B(G330), .C1(new_n934), .C2(new_n936), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n709), .A3(new_n968), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1157), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT116), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n742), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1164), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT116), .B1(new_n1169), .B2(new_n747), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1150), .A2(new_n1164), .A3(new_n1156), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n835), .A2(G128), .B1(new_n808), .B2(G132), .ZN(new_n1173));
  INV_X1    g0973(.A(G125), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n262), .C1(new_n1174), .C2(new_n813), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n1121), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT53), .B1(new_n825), .B2(new_n1121), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n406), .B2(new_n816), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT54), .B(G143), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1181), .A2(new_n806), .B1(new_n885), .B2(new_n822), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT117), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1179), .B(new_n1183), .C1(new_n211), .C2(new_n820), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n823), .A2(new_n322), .B1(new_n808), .B2(G116), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n568), .B2(new_n806), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n833), .A2(G294), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n835), .A2(G283), .B1(new_n839), .B2(G77), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n262), .B(new_n881), .C1(G87), .C2(new_n897), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1184), .A2(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1192), .A2(new_n878), .B1(new_n334), .B2(new_n875), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n804), .B(new_n1193), .C1(new_n1151), .C2(new_n854), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1157), .B2(new_n1051), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT118), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT118), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1131), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n1194), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1172), .A2(new_n1200), .ZN(G378));
  XNOR2_X1  g1001(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n708), .A2(new_n370), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n354), .A2(new_n904), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n708), .A2(new_n370), .A3(new_n1207), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1207), .B1(new_n708), .B2(new_n370), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n696), .B(new_n1208), .C1(new_n706), .C2(new_n707), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1204), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1203), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(new_n1210), .A3(new_n1205), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1204), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1202), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1219), .A2(G330), .A3(new_n941), .A4(new_n948), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n868), .B(new_n929), .C1(new_n934), .C2(new_n936), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n922), .B2(new_n921), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G330), .B(new_n948), .C1(new_n1222), .C2(KEYINPUT40), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1216), .A2(new_n1217), .A3(new_n1202), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1202), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1220), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n966), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n963), .A2(new_n1220), .A3(new_n1227), .A4(new_n965), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1131), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1226), .A2(new_n855), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n818), .A2(new_n1174), .B1(new_n816), .B2(new_n1121), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT119), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n807), .A2(G137), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G132), .A2(new_n823), .B1(new_n897), .B2(new_n1180), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n808), .A2(G128), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT59), .Z(new_n1239));
  AOI21_X1  g1039(.A(G41), .B1(new_n833), .B2(G124), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G33), .B1(new_n981), .B2(G159), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n820), .A2(new_n201), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G283), .B2(new_n833), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1083), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n1005), .A2(new_n806), .B1(new_n202), .B2(new_n816), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1245), .A2(G41), .A3(new_n262), .A4(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G97), .A2(new_n823), .B1(new_n835), .B2(G116), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n215), .C2(new_n890), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT58), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n211), .B1(new_n357), .B2(G41), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1242), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n843), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT120), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(G50), .B2(new_n875), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1232), .A2(new_n804), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1231), .A2(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n968), .A2(new_n709), .A3(new_n1163), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1166), .A2(new_n1260), .B1(new_n1230), .B2(new_n1229), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n742), .B1(new_n1261), .B2(KEYINPUT57), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n968), .A2(new_n709), .A3(new_n1163), .ZN(new_n1263));
  AND4_X1   g1063(.A1(new_n965), .A2(new_n963), .A3(new_n1220), .A4(new_n1227), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n965), .A2(new_n963), .B1(new_n1220), .B2(new_n1227), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1263), .A2(new_n1169), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT57), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1259), .B1(new_n1262), .B2(new_n1268), .ZN(G375));
  OAI22_X1  g1069(.A1(new_n890), .A2(new_n885), .B1(new_n818), .B2(new_n879), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n806), .A2(new_n1121), .B1(new_n816), .B2(new_n211), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT123), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n414), .B(new_n1243), .C1(G128), .C2(new_n833), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1272), .B(new_n1273), .C1(new_n406), .C2(new_n825), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1270), .B1(new_n1274), .B2(KEYINPUT124), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(KEYINPUT124), .B2(new_n1274), .C1(new_n822), .C2(new_n1181), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n813), .A2(new_n633), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n890), .A2(new_n830), .B1(new_n818), .B2(new_n891), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G116), .B2(new_n823), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n807), .A2(new_n322), .B1(new_n839), .B2(new_n335), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n414), .B1(new_n820), .B2(new_n337), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G97), .B2(new_n897), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1276), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n843), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(G68), .B2(new_n875), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n804), .B(new_n1286), .C1(new_n854), .C2(new_n1139), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1162), .B2(new_n1051), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1070), .B1(new_n1260), .B2(new_n1162), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1165), .ZN(G381));
  OR2_X1    g1090(.A1(new_n1231), .A2(new_n1258), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n747), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1166), .A2(new_n1260), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(KEYINPUT57), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1291), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1011), .B(new_n1135), .C1(new_n1050), .C2(new_n1071), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1105), .A2(new_n860), .A3(new_n803), .A4(new_n1108), .ZN(new_n1298));
  NOR4_X1   g1098(.A1(new_n1297), .A2(G384), .A3(G381), .A4(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1172), .A2(new_n1200), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .ZN(G407));
  NOR2_X1   g1101(.A1(new_n1299), .A2(new_n716), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1303));
  OAI21_X1  g1103(.A(G213), .B1(new_n1302), .B2(new_n1303), .ZN(G409));
  NAND2_X1  g1104(.A1(new_n716), .A2(G213), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1293), .A2(new_n1070), .A3(new_n1294), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1172), .A2(new_n1200), .A3(new_n1259), .A4(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1305), .B(new_n1307), .C1(new_n1296), .C2(new_n1300), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1263), .A2(KEYINPUT60), .A3(new_n1161), .A4(new_n1159), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1260), .B2(new_n1162), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n747), .B1(new_n1260), .B2(new_n1162), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1162), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(KEYINPUT125), .A3(new_n1263), .A4(KEYINPUT60), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1288), .ZN(new_n1318));
  INV_X1    g1118(.A(G384), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT126), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1317), .A2(G384), .A3(new_n1288), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1318), .A2(new_n1323), .A3(new_n1319), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1321), .A2(new_n1322), .A3(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT62), .B1(new_n1308), .B2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n716), .A2(G213), .A3(G2897), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1323), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1329));
  AOI211_X1 g1129(.A(KEYINPUT126), .B(G384), .C1(new_n1317), .C2(new_n1288), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1328), .B1(new_n1331), .B2(new_n1322), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1322), .ZN(new_n1333));
  NOR4_X1   g1133(.A1(new_n1329), .A2(new_n1330), .A3(new_n1333), .A4(new_n1327), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1295), .A3(new_n742), .ZN(new_n1336));
  AOI22_X1  g1136(.A1(new_n1336), .A2(new_n1259), .B1(new_n1200), .B2(new_n1172), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1307), .A2(new_n1305), .ZN(new_n1338));
  OAI22_X1  g1138(.A1(new_n1332), .A2(new_n1334), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT61), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1307), .A2(new_n1305), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G375), .A2(G378), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1329), .A2(new_n1330), .A3(new_n1333), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .A4(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1326), .A2(new_n1339), .A3(new_n1340), .A4(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G387), .A2(G390), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G393), .A2(G396), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1298), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1348), .A2(new_n1350), .A3(new_n1297), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1350), .B1(new_n1348), .B2(new_n1297), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1347), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1349), .A2(new_n1298), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1297), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1070), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1356), .B1(new_n1133), .B2(new_n1053), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1046), .B(new_n1049), .C1(new_n1357), .C2(new_n1051), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1135), .B1(new_n1358), .B2(new_n1011), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1354), .B1(new_n1355), .B2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1348), .A2(new_n1350), .A3(new_n1297), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1360), .A2(KEYINPUT127), .A3(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1353), .A2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1346), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1360), .A2(new_n1340), .A3(new_n1361), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1337), .A2(new_n1338), .A3(new_n1325), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1365), .B1(new_n1366), .B2(KEYINPUT63), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT63), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1331), .A2(new_n1322), .A3(new_n1328), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1368), .B1(new_n1371), .B2(new_n1308), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1367), .B1(new_n1372), .B2(new_n1366), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1364), .A2(new_n1373), .ZN(G405));
  AND3_X1   g1174(.A1(new_n1360), .A2(KEYINPUT127), .A3(new_n1361), .ZN(new_n1375));
  AOI21_X1  g1175(.A(KEYINPUT127), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1376));
  OAI211_X1 g1176(.A(new_n1303), .B(new_n1342), .C1(new_n1375), .C2(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1342), .A2(new_n1303), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1378), .A2(new_n1353), .A3(new_n1362), .ZN(new_n1379));
  AND3_X1   g1179(.A1(new_n1377), .A2(new_n1344), .A3(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1344), .B1(new_n1377), .B2(new_n1379), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1380), .A2(new_n1381), .ZN(G402));
endmodule


