//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G85gat), .Z(new_n204));
  XNOR2_X1  g003(.A(G1gat), .B(G29gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n210), .B2(KEYINPUT68), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT68), .B2(new_n210), .ZN(new_n212));
  XOR2_X1   g011(.A(G127gat), .B(G134gat), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G120gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(G113gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT69), .B(G113gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G120gat), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n218), .A2(KEYINPUT1), .A3(new_n213), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(G141gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(KEYINPUT70), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(KEYINPUT70), .B2(new_n223), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  OR2_X1    g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(KEYINPUT2), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n223), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(new_n222), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n226), .B(new_n227), .C1(new_n231), .C2(KEYINPUT2), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n220), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT73), .Z(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n234), .B2(new_n220), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT71), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(KEYINPUT4), .B2(new_n236), .ZN(new_n244));
  INV_X1    g043(.A(new_n220), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n239), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n244), .A2(KEYINPUT74), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT74), .B1(new_n244), .B2(new_n251), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT5), .B(new_n240), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  INV_X1    g054(.A(new_n235), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n236), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OR3_X1    g057(.A1(new_n258), .A2(KEYINPUT5), .A3(new_n239), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n209), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n203), .B1(new_n260), .B2(KEYINPUT6), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n203), .A3(KEYINPUT6), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n254), .A2(new_n209), .A3(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n259), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n208), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n260), .A2(KEYINPUT79), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  INV_X1    g075(.A(G218gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(KEYINPUT22), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G211gat), .B(G218gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n247), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT3), .B1(new_n281), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n234), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G22gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G78gat), .B(G106gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT31), .B(G50gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n288), .B(new_n289), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT28), .Z(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT67), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n306), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(KEYINPUT26), .B2(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n312), .B2(new_n314), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT23), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n319), .C1(new_n304), .C2(new_n305), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n311), .B1(new_n313), .B2(new_n303), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n323), .A2(new_n324), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n309), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(new_n220), .ZN(new_n331));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT64), .Z(new_n333));
  NOR2_X1   g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT34), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT34), .B1(new_n334), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(new_n333), .ZN(new_n339));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  OAI211_X1 g141(.A(new_n339), .B(new_n342), .C1(new_n334), .C2(KEYINPUT33), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT33), .ZN(new_n344));
  INV_X1    g143(.A(new_n342), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n331), .B(new_n333), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n336), .A2(new_n343), .A3(new_n337), .A4(new_n346), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n298), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n330), .A2(new_n282), .B1(G226gat), .B2(G233gat), .ZN(new_n352));
  AND2_X1   g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n330), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(new_n281), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n281), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n357), .B2(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n364), .A3(new_n362), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n202), .B1(new_n274), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n269), .A2(new_n266), .A3(new_n265), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n262), .A2(new_n371), .A3(new_n263), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n296), .B(new_n297), .ZN(new_n373));
  INV_X1    g172(.A(new_n350), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT36), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT36), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n350), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n298), .A2(new_n202), .A3(new_n350), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n372), .B(new_n368), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n361), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(KEYINPUT38), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT38), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n271), .A2(new_n272), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n258), .A2(new_n239), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(KEYINPUT39), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n237), .A2(new_n239), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT39), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n389), .B2(KEYINPUT78), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n209), .B(new_n390), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT40), .ZN(new_n396));
  INV_X1    g195(.A(new_n368), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n274), .A2(new_n387), .B1(new_n388), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n375), .ZN(new_n400));
  INV_X1    g199(.A(new_n377), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n373), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n370), .B(new_n380), .C1(new_n399), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G15gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n289), .ZN(new_n405));
  INV_X1    g204(.A(G1gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(G15gat), .A2(G22gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n409));
  AOI21_X1  g208(.A(G8gat), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n411));
  INV_X1    g210(.A(new_n407), .ZN(new_n412));
  NOR2_X1   g211(.A1(G15gat), .A2(G22gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n408), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n414), .B(new_n408), .C1(new_n409), .C2(G8gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G43gat), .B(G50gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n422));
  INV_X1    g221(.A(G29gat), .ZN(new_n423));
  INV_X1    g222(.A(G36gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G29gat), .A2(G36gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n427), .B2(new_n426), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT15), .B(new_n421), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G43gat), .B(G50gat), .Z(new_n433));
  INV_X1    g232(.A(KEYINPUT15), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n421), .A2(KEYINPUT15), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n425), .A2(new_n427), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n430), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT84), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n430), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n437), .B1(KEYINPUT15), .B2(new_n421), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n431), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n436), .B1(new_n446), .B2(new_n428), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n442), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n438), .A3(KEYINPUT17), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n418), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(KEYINPUT18), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n439), .ZN(new_n454));
  INV_X1    g253(.A(new_n440), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT84), .B1(new_n416), .B2(new_n417), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(KEYINPUT85), .A3(new_n441), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n420), .A2(new_n459), .A3(new_n439), .A4(new_n440), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n452), .B(KEYINPUT13), .Z(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n453), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n441), .A2(new_n450), .A3(new_n452), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT18), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n469));
  XNOR2_X1  g268(.A(G113gat), .B(G141gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G169gat), .B(G197gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT12), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n467), .A2(KEYINPUT86), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n465), .A2(new_n479), .A3(new_n466), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n478), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n474), .A3(new_n480), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n483), .A2(new_n463), .A3(KEYINPUT87), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n476), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT21), .ZN(new_n486));
  AND2_X1   g285(.A1(G71gat), .A2(G78gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G57gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(G64gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT88), .B(G57gat), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(G64gat), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n491), .A2(G71gat), .A3(G78gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(new_n487), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n455), .A2(new_n456), .B1(new_n486), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT91), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT19), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n501), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G127gat), .B(G155gat), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT20), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n504), .B(new_n506), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n486), .ZN(new_n508));
  XNOR2_X1  g307(.A(G183gat), .B(G211gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G231gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n507), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G99gat), .B(G106gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT93), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(KEYINPUT93), .A3(new_n521), .ZN(new_n524));
  NOR2_X1   g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT8), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n516), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n525), .B1(new_n531), .B2(new_n517), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n515), .A4(new_n528), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n448), .A2(new_n449), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n537), .C1(new_n454), .C2(new_n535), .ZN(new_n538));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT92), .ZN(new_n542));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT94), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n544), .B(KEYINPUT94), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n540), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n514), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G176gat), .B(G204gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT96), .ZN(new_n553));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT10), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n535), .A2(new_n557), .A3(new_n499), .ZN(new_n558));
  AND2_X1   g357(.A1(KEYINPUT88), .A2(G57gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT88), .A2(G57gat), .ZN(new_n560));
  OAI21_X1  g359(.A(G64gat), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n493), .B2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n498), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n493), .A2(G64gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT9), .B1(new_n564), .B2(new_n494), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n562), .A2(new_n563), .B1(new_n565), .B2(new_n489), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n534), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n535), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n534), .B(new_n530), .C1(new_n499), .C2(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n558), .B1(new_n571), .B2(new_n557), .ZN(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT97), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT98), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT10), .B1(new_n569), .B2(new_n570), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n577), .B(new_n574), .C1(new_n578), .C2(new_n558), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n571), .A2(new_n573), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n556), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n573), .B1(new_n578), .B2(new_n558), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n555), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND4_X1   g386(.A1(new_n403), .A2(new_n485), .A3(new_n551), .A4(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n372), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT99), .B(G1gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(G1324gat));
  XOR2_X1   g391(.A(KEYINPUT16), .B(G8gat), .Z(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n397), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT42), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT42), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n397), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n597), .B2(G8gat), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n594), .B2(new_n598), .ZN(G1325gat));
  AOI21_X1  g398(.A(G15gat), .B1(new_n588), .B2(new_n374), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n400), .A2(new_n401), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n404), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n588), .B2(new_n603), .ZN(G1326gat));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n298), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT43), .B(G22gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(G1327gat));
  INV_X1    g406(.A(new_n263), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n261), .ZN(new_n609));
  INV_X1    g408(.A(new_n267), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n269), .A2(new_n270), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n260), .A2(KEYINPUT79), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n369), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n380), .B1(new_n614), .B2(KEYINPUT35), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n387), .A2(new_n609), .A3(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n398), .A2(new_n388), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n402), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n550), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n485), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n513), .A2(new_n621), .A3(new_n586), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n623), .A2(G29gat), .A3(new_n372), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT45), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n403), .B2(new_n550), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n631), .B(new_n550), .C1(new_n615), .C2(new_n618), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n622), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(G29gat), .B1(new_n635), .B2(new_n372), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n626), .A2(KEYINPUT45), .A3(new_n627), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n630), .A2(new_n636), .A3(new_n637), .ZN(G1328gat));
  NOR3_X1   g437(.A1(new_n623), .A2(G36gat), .A3(new_n368), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT101), .B(KEYINPUT46), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(G36gat), .B1(new_n635), .B2(new_n368), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(G1329gat));
  INV_X1    g442(.A(new_n623), .ZN(new_n644));
  INV_X1    g443(.A(G43gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n374), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n635), .A2(new_n602), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(new_n645), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g448(.A(G50gat), .B1(new_n635), .B2(new_n373), .ZN(new_n650));
  INV_X1    g449(.A(G50gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n298), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g455(.A1(new_n514), .A2(new_n485), .A3(new_n550), .A4(new_n587), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n403), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n403), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n372), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n495), .ZN(G1332gat));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(KEYINPUT104), .A3(new_n661), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n397), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT49), .B(G64gat), .Z(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n668), .B2(new_n670), .ZN(G1333gat));
  NAND4_X1  g470(.A1(new_n666), .A2(G71gat), .A3(new_n601), .A4(new_n667), .ZN(new_n672));
  INV_X1    g471(.A(G71gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n662), .B2(new_n350), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT50), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT50), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(G1334gat));
  NAND3_X1  g478(.A1(new_n666), .A2(new_n298), .A3(new_n667), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT105), .B(G78gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1335gat));
  NOR2_X1   g481(.A1(new_n513), .A2(new_n485), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT51), .B1(new_n619), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT51), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n403), .A2(new_n686), .A3(new_n550), .A4(new_n683), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n685), .A2(new_n687), .A3(new_n586), .ZN(new_n688));
  AOI21_X1  g487(.A(G85gat), .B1(new_n688), .B2(new_n589), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n587), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n619), .A2(KEYINPUT44), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n633), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n589), .A2(G85gat), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n689), .B1(new_n693), .B2(new_n694), .ZN(G1336gat));
  OAI211_X1 g494(.A(new_n397), .B(new_n690), .C1(new_n632), .C2(new_n634), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G92gat), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT52), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G92gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n693), .B2(new_n397), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n368), .A2(G92gat), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n685), .A2(new_n687), .A3(new_n586), .A4(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT107), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n697), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n699), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n697), .A2(new_n698), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n705), .A2(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n708), .A2(new_n711), .ZN(G1337gat));
  AOI21_X1  g511(.A(G99gat), .B1(new_n688), .B2(new_n374), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n601), .A2(G99gat), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n693), .B2(new_n714), .ZN(G1338gat));
  INV_X1    g514(.A(KEYINPUT53), .ZN(new_n716));
  INV_X1    g515(.A(G106gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n688), .A2(new_n717), .A3(new_n298), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n693), .A2(new_n298), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI221_X1 g522(.A(new_n718), .B1(new_n719), .B2(new_n716), .C1(new_n717), .C2(new_n721), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1339gat));
  NAND2_X1  g524(.A1(new_n589), .A2(new_n368), .ZN(new_n726));
  INV_X1    g525(.A(new_n351), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n585), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n572), .A2(new_n575), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(KEYINPUT54), .A3(new_n583), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT54), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n580), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n735), .A3(new_n556), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT54), .B1(new_n576), .B2(new_n579), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n737), .B2(new_n555), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n732), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n729), .B1(new_n739), .B2(KEYINPUT55), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n735), .B1(new_n734), .B2(new_n556), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n555), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n731), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n740), .A2(new_n485), .A3(new_n745), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n482), .A2(new_n484), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n461), .B1(new_n458), .B2(new_n460), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n451), .A2(new_n452), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n473), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT110), .Z(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n586), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n550), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT55), .B(new_n731), .C1(new_n741), .C2(new_n742), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n745), .A2(new_n550), .A3(new_n585), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n747), .A2(new_n751), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n514), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n550), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n513), .A2(new_n621), .A3(new_n759), .A4(new_n587), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n728), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n621), .ZN(new_n763));
  MUX2_X1   g562(.A(G113gat), .B(new_n217), .S(new_n763), .Z(G1340gat));
  OAI21_X1  g563(.A(G120gat), .B1(new_n762), .B2(new_n587), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n586), .A2(new_n215), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n762), .B2(new_n767), .ZN(G1341gat));
  NOR2_X1   g567(.A1(new_n762), .A2(new_n514), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g569(.A1(new_n762), .A2(new_n759), .ZN(new_n771));
  INV_X1    g570(.A(G134gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(KEYINPUT56), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(KEYINPUT56), .B2(new_n774), .ZN(G1343gat));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n726), .A2(new_n601), .ZN(new_n778));
  INV_X1    g577(.A(new_n757), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n485), .B1(new_n739), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n754), .A2(new_n585), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n752), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n759), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n513), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n760), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT57), .B(new_n298), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT113), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n373), .B1(new_n758), .B2(new_n760), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(KEYINPUT57), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n778), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(new_n621), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G141gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n621), .A2(G141gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT114), .Z(new_n796));
  AOI21_X1  g595(.A(new_n777), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n799), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n777), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n792), .B2(G141gat), .ZN(new_n803));
  OR3_X1    g602(.A1(new_n797), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n797), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1344gat));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n756), .B1(new_n755), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n740), .A2(new_n745), .A3(KEYINPUT118), .A4(new_n550), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n513), .B1(new_n811), .B2(new_n784), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT119), .B1(new_n812), .B2(new_n786), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n809), .A2(new_n810), .B1(new_n759), .B2(new_n783), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n814), .B(new_n760), .C1(new_n815), .C2(new_n513), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n298), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(KEYINPUT120), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n789), .A2(KEYINPUT57), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n760), .B1(new_n815), .B2(new_n513), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n373), .B1(new_n822), .B2(KEYINPUT119), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n823), .B2(new_n816), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(KEYINPUT120), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n726), .A2(KEYINPUT117), .A3(new_n601), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n778), .A2(new_n828), .ZN(new_n829));
  OR4_X1    g628(.A1(new_n587), .A2(new_n826), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n807), .B1(new_n830), .B2(G148gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n791), .A2(new_n587), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(KEYINPUT59), .A3(new_n221), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n778), .A2(new_n789), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n586), .A2(new_n221), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n831), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(G1345gat));
  INV_X1    g635(.A(G155gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n791), .A2(new_n837), .A3(new_n514), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n778), .A2(new_n513), .A3(new_n789), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n791), .B2(new_n759), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n759), .A2(G162gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n834), .B2(new_n842), .ZN(G1347gat));
  AND2_X1   g642(.A1(new_n761), .A2(new_n372), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n727), .A2(new_n368), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n621), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(new_n304), .ZN(G1348gat));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n587), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT121), .B(G176gat), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(G1349gat));
  NOR2_X1   g650(.A1(new_n846), .A2(new_n514), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT122), .B1(new_n852), .B2(new_n299), .ZN(new_n853));
  INV_X1    g652(.A(G183gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n852), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g655(.A1(new_n844), .A2(new_n550), .A3(new_n845), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(G190gat), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT123), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(G190gat), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT61), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1351gat));
  OR2_X1    g661(.A1(new_n826), .A2(KEYINPUT124), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n826), .A2(KEYINPUT124), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n589), .A2(new_n601), .A3(new_n368), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G197gat), .B1(new_n866), .B2(new_n621), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n378), .A2(new_n397), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n844), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n621), .A2(G197gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(G1352gat));
  OAI21_X1  g670(.A(G204gat), .B1(new_n866), .B2(new_n587), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n869), .A2(G204gat), .A3(new_n587), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT62), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1353gat));
  NAND4_X1  g674(.A1(new_n844), .A2(new_n276), .A3(new_n513), .A4(new_n868), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n865), .A2(new_n513), .ZN(new_n878));
  INV_X1    g677(.A(new_n820), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n824), .B2(KEYINPUT120), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n817), .A2(new_n818), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT125), .B(new_n877), .C1(new_n884), .C2(new_n276), .ZN(new_n885));
  INV_X1    g684(.A(new_n878), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n821), .B2(new_n825), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(G211gat), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT125), .B1(new_n890), .B2(new_n877), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n876), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT126), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n894), .B(new_n876), .C1(new_n889), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1354gat));
  INV_X1    g695(.A(new_n866), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n550), .A2(G218gat), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT127), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n844), .A2(new_n550), .A3(new_n868), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n897), .A2(new_n899), .B1(new_n277), .B2(new_n900), .ZN(G1355gat));
endmodule


