//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n993, new_n994,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1058, new_n1059;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G134gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(G120gat), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  INV_X1    g015(.A(G120gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G113gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n215), .B2(new_n218), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n212), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT78), .ZN(new_n230));
  AND2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(KEYINPUT78), .A3(new_n224), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G141gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n242), .B2(G148gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n229), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n224), .ZN(new_n246));
  XOR2_X1   g045(.A(G141gat), .B(G148gat), .Z(new_n247));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n240), .A2(new_n241), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n238), .B1(new_n251), .B2(new_n237), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n214), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n254), .A2(new_n255), .A3(new_n217), .ZN(new_n256));
  INV_X1    g055(.A(new_n218), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(new_n219), .A3(new_n220), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(new_n212), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n203), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(new_n223), .B2(new_n244), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n253), .A2(new_n259), .A3(KEYINPUT4), .A4(new_n212), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n244), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n269), .B(new_n229), .C1(new_n236), .C2(new_n243), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n270), .A3(new_n223), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT79), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n266), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n264), .B1(new_n273), .B2(new_n263), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n266), .A2(new_n267), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n253), .B2(new_n269), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n268), .A3(new_n270), .A4(new_n223), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n275), .A2(new_n203), .A3(new_n262), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT0), .ZN(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G85gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n202), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n274), .B2(new_n279), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n284), .A3(new_n279), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT35), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301));
  INV_X1    g100(.A(G211gat), .ZN(new_n302));
  INV_X1    g101(.A(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n300), .A3(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n318), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n331), .A2(G169gat), .A3(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n314), .B1(new_n325), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n316), .A2(new_n317), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n319), .B1(new_n337), .B2(KEYINPUT24), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n322), .B(new_n336), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(KEYINPUT66), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(KEYINPUT23), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n314), .B1(new_n327), .B2(new_n329), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G183gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n349), .A3(new_n317), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT28), .A3(new_n317), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n319), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n357), .A3(new_n343), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n359), .A2(new_n328), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n335), .A2(new_n346), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n313), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n361), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n332), .B1(new_n327), .B2(new_n329), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT25), .B1(new_n367), .B2(new_n324), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n313), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n312), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n363), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT74), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n311), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n313), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n310), .A3(new_n371), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(KEYINPUT75), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n382), .B(new_n311), .C1(new_n372), .C2(new_n375), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n299), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n298), .B(KEYINPUT76), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n362), .A2(new_n313), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT74), .B1(new_n374), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n364), .A2(new_n312), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n310), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n383), .B(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT30), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n383), .B1(new_n390), .B2(new_n391), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT30), .B1(new_n395), .B2(new_n298), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n204), .A2(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n219), .A2(new_n220), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n258), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n369), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT64), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n335), .A2(new_n346), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n223), .A3(new_n365), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n408));
  XOR2_X1   g207(.A(G15gat), .B(G43gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT70), .ZN(new_n410));
  XOR2_X1   g209(.A(G71gat), .B(G99gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n407), .B2(KEYINPUT32), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n407), .A2(new_n413), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT71), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n404), .ZN(new_n423));
  INV_X1    g222(.A(new_n406), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n362), .A2(new_n223), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT34), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n423), .C1(new_n424), .C2(new_n425), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n417), .A2(new_n418), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT71), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n419), .ZN(new_n435));
  INV_X1    g234(.A(new_n430), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n416), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n363), .B1(new_n308), .B2(new_n309), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n244), .B1(new_n439), .B2(KEYINPUT3), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT82), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n310), .B1(new_n270), .B2(new_n373), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G228gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(new_n244), .C1(new_n439), .C2(KEYINPUT3), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n441), .A2(new_n443), .A3(new_n444), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n310), .A2(new_n377), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n253), .B1(new_n448), .B2(new_n269), .ZN(new_n449));
  OAI211_X1 g248(.A(G228gat), .B(G233gat), .C1(new_n449), .C2(new_n442), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n447), .B2(new_n450), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n438), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G78gat), .B(G106gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(G22gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n450), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  INV_X1    g258(.A(new_n438), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n452), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n457), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n457), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n453), .A2(new_n454), .A3(new_n438), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n460), .B1(new_n459), .B2(new_n452), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n431), .A2(new_n437), .A3(new_n462), .A4(new_n466), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n295), .A2(new_n398), .A3(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n291), .A2(KEYINPUT80), .A3(new_n287), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT80), .B1(new_n291), .B2(new_n287), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n469), .A2(new_n470), .A3(new_n289), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n288), .A2(new_n290), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n394), .B(new_n397), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT35), .B1(new_n473), .B2(new_n467), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n291), .A2(new_n287), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n291), .A2(KEYINPUT80), .A3(new_n287), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n286), .A3(new_n480), .ZN(new_n481));
  AND4_X1   g280(.A1(KEYINPUT81), .A2(new_n280), .A3(KEYINPUT6), .A4(new_n285), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT81), .B1(new_n289), .B2(KEYINPUT6), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n395), .A2(new_n298), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n392), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n396), .B1(new_n487), .B2(KEYINPUT30), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n436), .B1(new_n435), .B2(new_n416), .ZN(new_n489));
  AOI211_X1 g288(.A(new_n415), .B(new_n430), .C1(new_n434), .C2(new_n419), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n466), .A2(new_n462), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n485), .A2(new_n488), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n273), .A2(new_n263), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(KEYINPUT39), .C1(new_n263), .C2(new_n261), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n273), .A2(new_n497), .A3(new_n263), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n498), .A2(KEYINPUT84), .A3(new_n284), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT84), .B1(new_n498), .B2(new_n284), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n289), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n486), .B2(new_n392), .ZN(new_n505));
  OAI221_X1 g304(.A(new_n503), .B1(new_n502), .B2(new_n501), .C1(new_n505), .C2(new_n396), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n395), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n299), .B1(new_n395), .B2(new_n507), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n310), .B1(new_n372), .B2(new_n375), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n387), .B1(new_n313), .B2(new_n378), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n507), .B1(new_n513), .B2(new_n311), .ZN(new_n514));
  AOI211_X1 g313(.A(KEYINPUT38), .B(new_n385), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n508), .A2(new_n515), .A3(KEYINPUT85), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT85), .B1(new_n508), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n484), .A2(new_n486), .A3(new_n292), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n506), .B(new_n492), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n491), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n431), .A2(new_n437), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  NAND2_X1  g324(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n492), .B1(new_n485), .B2(new_n488), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n476), .A2(new_n494), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G43gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(G50gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT15), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G29gat), .ZN(new_n539));
  INV_X1    g338(.A(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT14), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n536), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G43gat), .B(G50gat), .Z(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n537), .B(KEYINPUT90), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n535), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT89), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n545), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  INV_X1    g355(.A(G1gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT16), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(G1gat), .B2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G8gat), .ZN(new_n561));
  INV_X1    g360(.A(G8gat), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n559), .B(new_n562), .C1(G1gat), .C2(new_n556), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n555), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n555), .A2(new_n564), .A3(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n564), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n535), .A2(new_n549), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n573), .A2(new_n548), .A3(new_n552), .A4(new_n553), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n574), .B2(new_n545), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n545), .B(new_n572), .C1(new_n550), .C2(new_n554), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n571), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n569), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n555), .A2(new_n564), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n569), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n570), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n579), .A2(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT88), .ZN(new_n587));
  XOR2_X1   g386(.A(G113gat), .B(G141gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n591), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT12), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT12), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n569), .A2(new_n578), .A3(KEYINPUT18), .A4(new_n570), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n585), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n585), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(G85gat), .B(G92gat), .C1(KEYINPUT98), .C2(KEYINPUT7), .ZN(new_n606));
  AND2_X1   g405(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n611));
  NAND2_X1  g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G99gat), .B(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(G99gat), .ZN(new_n615));
  INV_X1    g414(.A(G106gat), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT8), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n609), .A2(new_n613), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n612), .ZN(new_n620));
  INV_X1    g419(.A(new_n610), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n619), .B1(new_n622), .B2(new_n608), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n575), .B2(new_n577), .ZN(new_n625));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  INV_X1    g427(.A(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n555), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n631));
  INV_X1    g430(.A(G232gat), .ZN(new_n632));
  INV_X1    g431(.A(G233gat), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n628), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  AOI211_X1 g435(.A(KEYINPUT99), .B(new_n634), .C1(new_n629), .C2(new_n555), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n625), .B(new_n627), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n624), .B1(new_n574), .B2(new_n545), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT99), .B1(new_n640), .B2(new_n634), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n630), .A2(new_n628), .A3(new_n635), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n627), .B1(new_n643), .B2(new_n625), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n605), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n625), .B1(new_n636), .B2(new_n637), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n626), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n603), .B(new_n604), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n638), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G230gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n633), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n653));
  NAND2_X1  g452(.A1(G71gat), .A2(G78gat), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT9), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(G57gat), .A2(G64gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(G57gat), .A2(G64gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G71gat), .B(G78gat), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT93), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(G71gat), .B2(G78gat), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n659), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n653), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G57gat), .B(G64gat), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(KEYINPUT94), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n665), .A2(new_n672), .A3(new_n624), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n618), .A2(new_n623), .A3(new_n670), .A4(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n665), .A2(new_n672), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT95), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n672), .A3(KEYINPUT95), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n624), .A2(new_n676), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n652), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n652), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(G120gat), .B(G148gat), .Z(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n687), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(G183gat), .B(G211gat), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT21), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G127gat), .B(G155gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n696), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n702), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n700), .A3(new_n695), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n707));
  NAND2_X1  g506(.A1(G231gat), .A2(G233gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n680), .A2(KEYINPUT21), .A3(new_n681), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n571), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n710), .B2(new_n571), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  INV_X1    g515(.A(new_n709), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n706), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n706), .B1(new_n715), .B2(new_n718), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n650), .B(new_n694), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n531), .A2(new_n600), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n485), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G1gat), .ZN(G1324gat));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726));
  INV_X1    g525(.A(new_n722), .ZN(new_n727));
  OAI21_X1  g526(.A(G8gat), .B1(new_n727), .B2(new_n488), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G8gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n722), .A2(new_n398), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n726), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n731), .A2(new_n726), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n732), .A2(KEYINPUT104), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1325gat));
  INV_X1    g535(.A(new_n528), .ZN(new_n737));
  OAI21_X1  g536(.A(G15gat), .B1(new_n727), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n524), .A2(G15gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n727), .B2(new_n739), .ZN(G1326gat));
  INV_X1    g539(.A(new_n492), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT43), .B(G22gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1327gat));
  NAND2_X1  g543(.A1(new_n715), .A2(new_n718), .ZN(new_n745));
  INV_X1    g544(.A(new_n706), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n706), .A2(new_n715), .A3(new_n718), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n687), .B(new_n692), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n598), .A2(new_n599), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n531), .A2(new_n650), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n539), .A3(new_n723), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT45), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n531), .B2(new_n650), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n645), .A2(new_n649), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n493), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT86), .B1(new_n493), .B2(KEYINPUT35), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(new_n761), .A3(new_n468), .ZN(new_n762));
  INV_X1    g561(.A(new_n529), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n520), .A2(new_n737), .A3(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(KEYINPUT44), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n753), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(new_n723), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n756), .B1(new_n769), .B2(new_n539), .ZN(G1328gat));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n540), .A3(new_n398), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT46), .Z(new_n772));
  AND2_X1   g571(.A1(new_n768), .A2(new_n398), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n540), .ZN(G1329gat));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n528), .A3(new_n765), .A4(new_n767), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G43gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT105), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n778), .A3(G43gat), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n524), .A2(G43gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n754), .A2(new_n780), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n776), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n784), .A2(new_n783), .A3(new_n776), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n782), .A2(KEYINPUT47), .B1(new_n785), .B2(new_n786), .ZN(G1330gat));
  NAND4_X1  g586(.A1(new_n758), .A2(new_n741), .A3(new_n765), .A4(new_n767), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G50gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n474), .A2(new_n475), .ZN(new_n790));
  INV_X1    g589(.A(new_n468), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n494), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n530), .A2(new_n520), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n492), .A2(G50gat), .A3(new_n650), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n794), .A2(new_n752), .A3(new_n751), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT48), .B1(new_n796), .B2(KEYINPUT107), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1331gat));
  AOI21_X1  g598(.A(new_n759), .B1(new_n747), .B2(new_n748), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n800), .A2(new_n600), .A3(new_n750), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n723), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g604(.A1(new_n802), .A2(new_n488), .ZN(new_n806));
  NOR2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  AND2_X1   g606(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n806), .B2(new_n807), .ZN(G1333gat));
  NOR3_X1   g609(.A1(new_n802), .A2(G71gat), .A3(new_n524), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n803), .A2(new_n528), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(G71gat), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g613(.A1(new_n803), .A2(new_n741), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(G78gat), .ZN(G1335gat));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n752), .A2(new_n749), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n650), .B1(new_n792), .B2(new_n793), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n818), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n820), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n822), .B2(new_n818), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT108), .B1(new_n531), .B2(new_n650), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n485), .A2(G85gat), .A3(new_n694), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n825), .A2(new_n694), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n766), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G85gat), .B1(new_n833), .B2(new_n485), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1336gat));
  NAND3_X1  g634(.A1(new_n766), .A2(new_n398), .A3(new_n832), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(new_n836), .B2(G92gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n488), .A2(G92gat), .A3(new_n694), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g639(.A(KEYINPUT109), .B(new_n817), .C1(new_n826), .C2(new_n827), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n827), .A2(new_n820), .A3(new_n819), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT51), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(new_n838), .B1(G92gat), .B2(new_n836), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n840), .B1(new_n846), .B2(new_n847), .ZN(G1337gat));
  NAND4_X1  g647(.A1(new_n829), .A2(new_n615), .A3(new_n491), .A4(new_n750), .ZN(new_n849));
  OAI21_X1  g648(.A(G99gat), .B1(new_n833), .B2(new_n737), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1338gat));
  NOR3_X1   g650(.A1(new_n492), .A2(G106gat), .A3(new_n694), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n841), .A2(new_n844), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n758), .A2(new_n741), .A3(new_n765), .A4(new_n832), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(G106gat), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n853), .B1(new_n824), .B2(new_n828), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT110), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AND4_X1   g661(.A1(KEYINPUT51), .A2(new_n827), .A3(new_n820), .A4(new_n819), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT51), .B1(new_n826), .B2(new_n827), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n855), .B2(G106gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n858), .A2(new_n869), .ZN(G1339gat));
  NAND3_X1  g669(.A1(new_n800), .A2(new_n600), .A3(new_n694), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT10), .B1(new_n673), .B2(new_n674), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n685), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n677), .A2(new_n683), .A3(new_n652), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n692), .B1(new_n684), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT55), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n687), .A2(new_n692), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT55), .B1(new_n876), .B2(new_n878), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT111), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n585), .A2(new_n596), .A3(new_n597), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n592), .A2(new_n593), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n582), .A2(new_n584), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n570), .B1(new_n569), .B2(new_n578), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n650), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT55), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n677), .A2(new_n683), .A3(new_n652), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(new_n684), .A3(new_n877), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n877), .B(new_n685), .C1(new_n872), .C2(new_n873), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n693), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n891), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT111), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n880), .A4(new_n879), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n883), .A2(new_n890), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n752), .A3(new_n898), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n750), .A2(new_n884), .A3(new_n888), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n902), .B2(new_n650), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n871), .B1(new_n903), .B2(new_n749), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(new_n492), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n723), .A2(new_n488), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n524), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G113gat), .B1(new_n909), .B2(new_n600), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n904), .A2(new_n723), .ZN(new_n911));
  AND4_X1   g710(.A1(new_n488), .A2(new_n911), .A3(new_n492), .A4(new_n491), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(new_n213), .A3(new_n214), .A4(new_n752), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(G1340gat));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n217), .A3(new_n750), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT112), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n908), .A2(new_n750), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G120gat), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT112), .B(new_n217), .C1(new_n908), .C2(new_n750), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT113), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n922), .B(new_n915), .C1(new_n918), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1341gat));
  INV_X1    g723(.A(new_n749), .ZN(new_n925));
  OAI21_X1  g724(.A(G127gat), .B1(new_n909), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n912), .A2(new_n209), .A3(new_n749), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1342gat));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n207), .A3(new_n759), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n930));
  OAI21_X1  g729(.A(G134gat), .B1(new_n909), .B2(new_n650), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G1343gat));
  NOR3_X1   g732(.A1(new_n528), .A2(new_n398), .A3(new_n492), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n911), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(G141gat), .A3(new_n600), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(KEYINPUT58), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n528), .A2(new_n906), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT114), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n896), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n882), .A2(KEYINPUT114), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n880), .B(new_n879), .C1(new_n598), .C2(new_n599), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n901), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(new_n650), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n925), .B1(new_n946), .B2(new_n899), .ZN(new_n947));
  AOI211_X1 g746(.A(new_n939), .B(new_n492), .C1(new_n947), .C2(new_n871), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT57), .B1(new_n904), .B2(new_n741), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n938), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n251), .B1(new_n950), .B2(new_n600), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n937), .A2(KEYINPUT116), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT116), .B1(new_n937), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(KEYINPUT115), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT115), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(new_n938), .C1(new_n948), .C2(new_n949), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n752), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n936), .B1(new_n957), .B2(new_n251), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT58), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n952), .A2(new_n953), .B1(new_n958), .B2(new_n959), .ZN(G1344gat));
  NAND2_X1  g759(.A1(new_n938), .A2(new_n750), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n492), .A2(new_n939), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n904), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT117), .B1(new_n721), .B2(new_n752), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n800), .A2(new_n965), .A3(new_n600), .A4(new_n694), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n896), .A2(new_n759), .A3(new_n880), .A4(new_n879), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT118), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n889), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n881), .A2(new_n882), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(KEYINPUT118), .A3(new_n759), .ZN(new_n972));
  AOI22_X1  g771(.A1(new_n945), .A2(new_n650), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n967), .B1(new_n973), .B2(new_n749), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT57), .B1(new_n974), .B2(new_n741), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n963), .B1(new_n975), .B2(KEYINPUT119), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT119), .ZN(new_n978));
  AOI211_X1 g777(.A(new_n978), .B(KEYINPUT57), .C1(new_n974), .C2(new_n741), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n961), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT59), .B1(new_n981), .B2(new_n237), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n954), .A2(new_n956), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n983), .A2(new_n694), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n237), .A2(KEYINPUT59), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(new_n935), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(new_n237), .A3(new_n750), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(G1345gat));
  OAI21_X1  g788(.A(G155gat), .B1(new_n983), .B2(new_n925), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n225), .A3(new_n749), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1346gat));
  OAI21_X1  g791(.A(G162gat), .B1(new_n983), .B2(new_n650), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n987), .A2(new_n226), .A3(new_n759), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1347gat));
  NAND2_X1  g794(.A1(new_n904), .A2(new_n485), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n996), .A2(new_n488), .A3(new_n467), .ZN(new_n997));
  INV_X1    g796(.A(G169gat), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n998), .A3(new_n752), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT121), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n398), .A2(new_n485), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n1001), .A2(new_n524), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n905), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT120), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT120), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n905), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(new_n752), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1000), .B1(new_n1009), .B2(G169gat), .ZN(new_n1010));
  AOI211_X1 g809(.A(KEYINPUT121), .B(new_n998), .C1(new_n1008), .C2(new_n752), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n999), .B1(new_n1010), .B2(new_n1011), .ZN(G1348gat));
  NAND2_X1  g811(.A1(new_n750), .A2(G176gat), .ZN(new_n1013));
  OR3_X1    g812(.A1(new_n1007), .A2(KEYINPUT123), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g813(.A(G176gat), .B1(new_n997), .B2(new_n750), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT122), .ZN(new_n1016));
  OAI21_X1  g815(.A(KEYINPUT123), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1017));
  AND3_X1   g816(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(G1349gat));
  NAND3_X1  g817(.A1(new_n997), .A2(new_n353), .A3(new_n749), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1007), .A2(new_n925), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1019), .B1(new_n1020), .B2(new_n316), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1021), .A2(KEYINPUT60), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT60), .ZN(new_n1023));
  OAI211_X1 g822(.A(new_n1023), .B(new_n1019), .C1(new_n1020), .C2(new_n316), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1022), .A2(new_n1024), .ZN(G1350gat));
  NAND3_X1  g824(.A1(new_n1004), .A2(new_n759), .A3(new_n1006), .ZN(new_n1026));
  AOI21_X1  g825(.A(KEYINPUT124), .B1(new_n1026), .B2(G190gat), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT61), .ZN(new_n1028));
  NOR2_X1   g827(.A1(new_n650), .A2(G190gat), .ZN(new_n1029));
  AOI22_X1  g828(.A1(new_n1027), .A2(new_n1028), .B1(new_n997), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1026), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(G1351gat));
  NOR4_X1   g832(.A1(new_n996), .A2(new_n488), .A3(new_n492), .A4(new_n528), .ZN(new_n1034));
  AOI21_X1  g833(.A(G197gat), .B1(new_n1034), .B2(new_n752), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n977), .A2(new_n980), .ZN(new_n1036));
  NOR2_X1   g835(.A1(new_n528), .A2(new_n1001), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g837(.A(new_n1038), .ZN(new_n1039));
  AND2_X1   g838(.A1(new_n752), .A2(G197gat), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(G1352gat));
  XOR2_X1   g840(.A(KEYINPUT125), .B(G204gat), .Z(new_n1042));
  AOI21_X1  g841(.A(new_n1042), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1034), .A2(new_n750), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g843(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1045));
  XNOR2_X1  g844(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  OAI21_X1  g845(.A(new_n1042), .B1(new_n1038), .B2(new_n694), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(new_n1047), .ZN(G1353gat));
  NAND3_X1  g847(.A1(new_n1034), .A2(new_n302), .A3(new_n749), .ZN(new_n1049));
  OAI211_X1 g848(.A(new_n749), .B(new_n1037), .C1(new_n976), .C2(new_n979), .ZN(new_n1050));
  AND3_X1   g849(.A1(new_n1050), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1051));
  AOI21_X1  g850(.A(KEYINPUT63), .B1(new_n1050), .B2(G211gat), .ZN(new_n1052));
  OAI21_X1  g851(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1054));
  INV_X1    g853(.A(KEYINPUT127), .ZN(new_n1055));
  OAI211_X1 g854(.A(new_n1055), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g855(.A1(new_n1054), .A2(new_n1056), .ZN(G1354gat));
  OAI21_X1  g856(.A(G218gat), .B1(new_n1038), .B2(new_n650), .ZN(new_n1058));
  NAND3_X1  g857(.A1(new_n1034), .A2(new_n303), .A3(new_n759), .ZN(new_n1059));
  NAND2_X1  g858(.A1(new_n1058), .A2(new_n1059), .ZN(G1355gat));
endmodule


