//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(G226), .B(G232), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G68), .B(G77), .Z(new_n233));
  XOR2_X1   g0033(.A(G50), .B(G58), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G351));
  NAND3_X1  g0039(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n204), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  OAI221_X1 g0050(.A(new_n245), .B1(new_n246), .B2(new_n247), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n212), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n241), .A2(new_n253), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n203), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G68), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n244), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT11), .B1(new_n251), .B2(new_n253), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT14), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n266), .A3(G274), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G238), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n267), .B2(new_n269), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G226), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G232), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G97), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n281), .A2(KEYINPUT68), .A3(new_n282), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n212), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT13), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n273), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n273), .B2(new_n289), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n261), .B(G169), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n286), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT68), .B1(new_n281), .B2(new_n282), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n294), .A2(new_n295), .A3(new_n266), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n267), .A2(new_n269), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT69), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT13), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n273), .A2(new_n289), .A3(new_n290), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G179), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n302), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n261), .B1(new_n305), .B2(G169), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT70), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(G169), .B1(new_n291), .B2(new_n292), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT70), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n309), .A2(new_n310), .A3(new_n303), .A4(new_n293), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n260), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n305), .A2(G200), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n301), .A2(G190), .A3(new_n302), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n260), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT3), .B(G33), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(G222), .A3(new_n275), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(G223), .A3(G1698), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n320), .C1(new_n247), .C2(new_n318), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n288), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n266), .A2(new_n268), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G274), .ZN(new_n325));
  AND2_X1   g0125(.A1(G1), .A2(G13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n265), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n324), .A2(G226), .B1(new_n264), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n256), .A2(G50), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT66), .ZN(new_n332));
  INV_X1    g0132(.A(new_n255), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n332), .A2(new_n333), .B1(G50), .B2(new_n240), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  INV_X1    g0135(.A(G150), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n246), .B1(new_n336), .B2(new_n249), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT65), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G50), .A2(G58), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n204), .B1(new_n340), .B2(new_n242), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n337), .B2(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n334), .B1(new_n343), .B2(new_n253), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n330), .B(new_n344), .C1(new_n345), .C2(new_n329), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n329), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G200), .B2(new_n329), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n344), .A2(KEYINPUT9), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n344), .A2(KEYINPUT9), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT10), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n349), .A2(new_n354), .A3(new_n350), .A4(new_n351), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n346), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT3), .ZN(new_n358));
  INV_X1    g0158(.A(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n204), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n361), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n242), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G58), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n242), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G58), .A2(G68), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n248), .A2(G159), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n357), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n253), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n364), .A2(new_n365), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n372), .B1(new_n377), .B2(G68), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n378), .B2(KEYINPUT16), .ZN(new_n379));
  OAI211_X1 g0179(.A(KEYINPUT71), .B(new_n357), .C1(new_n366), .C2(new_n372), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n335), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n256), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n333), .A2(new_n383), .B1(new_n240), .B2(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n274), .A2(G1698), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n318), .B(new_n387), .C1(G223), .C2(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n266), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n267), .B1(new_n277), .B2(new_n323), .ZN(new_n391));
  OAI21_X1  g0191(.A(G169), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n288), .ZN(new_n394));
  INV_X1    g0194(.A(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n386), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT18), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n390), .A2(new_n391), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n381), .A2(new_n385), .B1(new_n392), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n347), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G200), .B2(new_n401), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n381), .A2(new_n407), .A3(new_n385), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n381), .A2(new_n407), .A3(KEYINPUT17), .A4(new_n385), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n400), .A2(new_n405), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G20), .A2(G77), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n414), .B1(new_n335), .B2(new_n249), .C1(new_n246), .C2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n253), .B1(new_n247), .B2(new_n241), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n256), .A2(G77), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT67), .B1(new_n333), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT67), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n255), .A2(new_n420), .A3(G77), .A4(new_n256), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n288), .B1(new_n318), .B2(G107), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n277), .A2(new_n275), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G238), .B2(new_n275), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n318), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G244), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n267), .B1(new_n428), .B2(new_n323), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n345), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n318), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n288), .C1(G107), .C2(new_n318), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n324), .A2(G244), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n397), .A3(new_n267), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n423), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(G200), .B1(new_n427), .B2(new_n429), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(G190), .A3(new_n267), .A4(new_n433), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n417), .A4(new_n422), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n317), .A2(new_n356), .A3(new_n413), .A4(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT78), .B(KEYINPUT21), .Z(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n241), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n376), .B(new_n240), .C1(G1), .C2(new_n359), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n442), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n204), .C1(G33), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n442), .A2(G20), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n253), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n253), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT20), .B(new_n448), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT72), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n263), .A2(G1), .ZN(new_n459));
  AND2_X1   g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(G274), .B1(new_n287), .B2(new_n212), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT5), .B(G41), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n327), .A2(KEYINPUT72), .A3(new_n465), .A4(new_n459), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n275), .A2(G264), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G257), .A2(G1698), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n468), .A2(new_n469), .B1(new_n279), .B2(new_n280), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n288), .C1(G303), .C2(new_n318), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n462), .A2(G270), .A3(new_n266), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n441), .B1(new_n457), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT79), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n477), .B(new_n441), .C1(new_n457), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n464), .A2(new_n466), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(G179), .A3(new_n472), .A4(new_n471), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n253), .A2(new_n450), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n253), .A2(new_n449), .A3(new_n450), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT20), .B1(new_n486), .B2(new_n448), .ZN(new_n487));
  INV_X1    g0287(.A(new_n456), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(KEYINPUT77), .B(new_n482), .C1(new_n489), .C2(new_n445), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT77), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n457), .B2(new_n481), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n457), .A2(new_n474), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n490), .A2(new_n492), .B1(new_n493), .B2(KEYINPUT21), .ZN(new_n494));
  OAI211_X1 g0294(.A(G257), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT81), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n318), .A2(KEYINPUT81), .A3(G257), .A4(G1698), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n318), .A2(G250), .A3(new_n275), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G294), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n288), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n465), .A2(new_n459), .B1(new_n326), .B2(new_n265), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G264), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n502), .A2(new_n504), .A3(new_n480), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n503), .B2(G264), .ZN(new_n507));
  AND4_X1   g0307(.A1(new_n506), .A2(new_n462), .A3(G264), .A4(new_n266), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n502), .A3(new_n480), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n505), .A2(new_n345), .B1(new_n510), .B2(new_n397), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  INV_X1    g0313(.A(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(G20), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n512), .A2(new_n515), .A3(new_n516), .A4(KEYINPUT80), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n204), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n318), .A2(new_n524), .A3(new_n204), .A4(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n521), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n253), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n240), .A2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT25), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n444), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G107), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n511), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n479), .A2(new_n494), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n480), .A2(new_n472), .A3(new_n471), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n539), .A2(new_n347), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(G200), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n457), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(G244), .C1(new_n280), .C2(new_n279), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n428), .B1(new_n360), .B2(new_n361), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n446), .C1(new_n546), .C2(KEYINPUT4), .ZN(new_n547));
  OAI21_X1  g0347(.A(G250), .B1(new_n279), .B2(new_n280), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n275), .B1(new_n548), .B2(KEYINPUT4), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n288), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n464), .A2(new_n466), .B1(new_n503), .B2(G257), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(G179), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n241), .A2(new_n447), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n444), .B2(new_n447), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n557), .A2(new_n447), .A3(G107), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n514), .B1(new_n364), .B2(new_n365), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n555), .B1(new_n565), .B2(new_n253), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n553), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT73), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n550), .A2(new_n568), .A3(new_n551), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n550), .B2(new_n551), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n345), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n552), .A2(KEYINPUT73), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n550), .A2(new_n568), .A3(new_n551), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(G190), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n559), .B1(new_n557), .B2(new_n556), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n576), .A2(new_n204), .B1(new_n247), .B2(new_n249), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n253), .B1(new_n577), .B2(new_n563), .ZN(new_n578));
  INV_X1    g0378(.A(new_n555), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G200), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n550), .B2(new_n551), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n572), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n204), .B1(new_n282), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  INV_X1    g0388(.A(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n204), .B(G68), .C1(new_n279), .C2(new_n280), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n586), .B1(new_n246), .B2(new_n447), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n253), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n415), .A2(new_n241), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT75), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n415), .B2(new_n444), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n266), .B1(G250), .B2(new_n459), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n263), .A2(G1), .A3(G274), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G238), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT74), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n318), .A2(new_n607), .A3(G244), .A4(G1698), .ZN(new_n608));
  OAI211_X1 g0408(.A(G244), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT74), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n603), .B1(new_n611), .B2(new_n266), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n345), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n608), .ZN(new_n614));
  INV_X1    g0414(.A(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n602), .B1(new_n616), .B2(new_n288), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n397), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n599), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n595), .A2(new_n596), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT75), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n596), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n612), .A2(G200), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n534), .A2(G87), .ZN(new_n626));
  OAI211_X1 g0426(.A(G190), .B(new_n603), .C1(new_n611), .C2(new_n266), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n505), .A2(new_n347), .B1(new_n510), .B2(new_n581), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n619), .B(new_n628), .C1(new_n629), .C2(new_n536), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n585), .A2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n440), .A2(new_n538), .A3(new_n542), .A4(new_n631), .ZN(G372));
  XNOR2_X1  g0432(.A(new_n403), .B(KEYINPUT18), .ZN(new_n633));
  INV_X1    g0433(.A(new_n435), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n312), .B1(new_n315), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n410), .A2(new_n411), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n353), .A2(new_n355), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n346), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n619), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n619), .A2(new_n628), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n580), .B1(G179), .B2(new_n552), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n573), .A2(new_n574), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n345), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(KEYINPUT26), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n619), .A2(new_n628), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n572), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n640), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n479), .A2(new_n494), .A3(new_n537), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n631), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n440), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n639), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(new_n537), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G343), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n509), .A2(new_n480), .A3(new_n502), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n502), .A2(new_n504), .A3(new_n480), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n663), .A2(G200), .B1(G190), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n530), .A3(new_n535), .ZN(new_n666));
  INV_X1    g0466(.A(new_n661), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n536), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n662), .B1(new_n669), .B2(new_n655), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n479), .A2(new_n494), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n661), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n662), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n457), .A2(new_n661), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n671), .B(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n542), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n674), .B1(new_n678), .B2(new_n670), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n590), .A2(G116), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n207), .A2(new_n262), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT84), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(new_n210), .B2(new_n683), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n685), .B2(new_n684), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT28), .Z(new_n688));
  AOI22_X1  g0488(.A1(new_n567), .A2(new_n571), .B1(new_n575), .B2(new_n583), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n641), .A2(new_n689), .A3(new_n666), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT87), .B1(new_n538), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT87), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n631), .A2(new_n692), .A3(new_n650), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n649), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(KEYINPUT29), .A3(new_n661), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT88), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n694), .A2(KEYINPUT88), .A3(KEYINPUT29), .A4(new_n661), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n667), .B1(new_n649), .B2(new_n651), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT85), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n482), .A2(new_n617), .A3(new_n502), .A4(new_n509), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n643), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n569), .A2(new_n570), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n509), .A2(new_n502), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n707), .A2(new_n612), .A3(new_n481), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n708), .A3(KEYINPUT30), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n539), .A2(new_n397), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n510), .A3(new_n552), .A4(new_n612), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n712), .B2(new_n667), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n702), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n667), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT85), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(KEYINPUT86), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n631), .A2(new_n538), .A3(new_n542), .A4(new_n661), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT86), .B1(new_n715), .B2(new_n719), .ZN(new_n723));
  OAI21_X1  g0523(.A(G330), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n701), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n688), .B1(new_n725), .B2(G1), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT89), .ZN(G364));
  INV_X1    g0527(.A(new_n683), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n204), .A2(G13), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n203), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n207), .A2(new_n318), .ZN(new_n734));
  INV_X1    g0534(.A(G355), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n735), .B1(G116), .B2(new_n207), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n235), .A2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n318), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n207), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n263), .B2(new_n211), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n736), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT90), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n212), .B1(G20), .B2(new_n345), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n733), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n746), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n204), .A2(new_n397), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n347), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G317), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT33), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n753), .A2(KEYINPUT33), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(G190), .A3(new_n581), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT94), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT93), .B(G326), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n761), .B(new_n762), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n347), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n204), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n204), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n772), .A2(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n318), .B1(new_n780), .B2(G329), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n750), .A2(new_n778), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n774), .A2(new_n347), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT92), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n777), .B(new_n784), .C1(G283), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n589), .B2(new_n775), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n318), .B1(new_n783), .B2(new_n247), .C1(new_n367), .C2(new_n758), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n751), .A2(new_n242), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n772), .A2(new_n447), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n768), .A2(G50), .B1(new_n790), .B2(G107), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n770), .A2(new_n791), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n745), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n748), .B1(new_n749), .B2(new_n801), .C1(new_n677), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n678), .A2(new_n733), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n677), .A2(G330), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n746), .A2(new_n743), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n733), .B1(new_n247), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n423), .A2(new_n667), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n438), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n435), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT99), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n423), .A2(new_n430), .A3(new_n434), .A4(new_n661), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n738), .B1(new_n780), .B2(G132), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n790), .A2(G68), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n250), .B2(new_n775), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT97), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n818), .B1(new_n367), .B2(new_n772), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n826));
  INV_X1    g0626(.A(new_n758), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT95), .B(G143), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n783), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n827), .A2(new_n829), .B1(new_n830), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n336), .B2(new_n751), .C1(new_n767), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT96), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT34), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n825), .A2(new_n826), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n789), .A2(new_n589), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G303), .B2(new_n768), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n783), .A2(new_n442), .B1(new_n779), .B2(new_n782), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n318), .B(new_n839), .C1(G294), .C2(new_n827), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n775), .A2(new_n514), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n841), .B(new_n798), .C1(G283), .C2(new_n752), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n808), .B1(new_n744), .B2(new_n817), .C1(new_n844), .C2(new_n749), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n699), .B(new_n817), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n724), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT101), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n732), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n724), .A2(new_n846), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n850), .B2(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n213), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n211), .B(G77), .C1(new_n367), .C2(new_n242), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n250), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n203), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n652), .A2(new_n661), .A3(new_n817), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n813), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n377), .A2(G68), .ZN(new_n865));
  INV_X1    g0665(.A(new_n372), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(KEYINPUT16), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n867), .A2(new_n253), .A3(new_n373), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(new_n384), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n660), .ZN(new_n870));
  INV_X1    g0670(.A(new_n636), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n633), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n386), .A2(new_n660), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n399), .A2(new_n873), .A3(new_n874), .A4(new_n408), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n868), .A2(new_n384), .B1(new_n398), .B2(new_n660), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n408), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n864), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n879), .C1(new_n413), .C2(new_n870), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n307), .A2(new_n311), .ZN(new_n884));
  INV_X1    g0684(.A(new_n260), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n260), .A2(new_n661), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n315), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n312), .B2(new_n316), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n863), .A2(new_n883), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n633), .B2(new_n660), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n381), .A2(new_n407), .A3(new_n385), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n659), .B1(new_n381), .B2(new_n385), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n895), .A2(new_n403), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT103), .B1(new_n897), .B2(new_n874), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n399), .A2(new_n873), .A3(new_n408), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT103), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT37), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n875), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n412), .A2(new_n896), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n870), .ZN(new_n905));
  AOI221_X4 g0705(.A(new_n864), .B1(new_n875), .B2(new_n878), .C1(new_n412), .C2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n894), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n312), .A2(new_n911), .A3(new_n661), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n312), .B2(new_n661), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n893), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n697), .A2(new_n440), .A3(new_n698), .A4(new_n700), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n639), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n721), .A2(new_n718), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n440), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT104), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n902), .A2(new_n903), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n906), .B1(new_n925), .B2(new_n864), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n888), .B1(new_n886), .B2(new_n315), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n312), .A2(new_n316), .A3(new_n887), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n922), .B(new_n817), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT40), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT40), .B1(new_n881), .B2(new_n882), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n816), .B1(new_n889), .B2(new_n890), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n922), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n924), .A2(new_n934), .ZN(new_n936));
  INV_X1    g0736(.A(G330), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n920), .A2(new_n938), .B1(new_n203), .B2(new_n729), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n920), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n861), .B1(new_n939), .B2(new_n940), .ZN(G367));
  OAI21_X1  g0741(.A(new_n689), .B1(new_n566), .B2(new_n661), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n644), .A2(new_n667), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT105), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n655), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n667), .B1(new_n947), .B2(new_n572), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n670), .A2(new_n672), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n944), .ZN(new_n951));
  XOR2_X1   g0751(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(KEYINPUT107), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT107), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n951), .B(new_n952), .Z(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n948), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n661), .B1(new_n624), .B2(new_n626), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n640), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n647), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT108), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n954), .A2(new_n957), .A3(new_n964), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n678), .A2(new_n670), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n946), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n954), .A2(new_n957), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n960), .B(KEYINPUT43), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n966), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n969), .B1(new_n966), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n944), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n673), .A2(KEYINPUT109), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT109), .B1(new_n673), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n673), .A2(new_n976), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT44), .Z(new_n983));
  NAND3_X1  g0783(.A1(new_n977), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n967), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n678), .A2(KEYINPUT110), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n670), .B(new_n672), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n725), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n725), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n683), .B(KEYINPUT41), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n730), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n975), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n747), .B1(new_n207), .B2(new_n415), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n231), .A2(new_n207), .A3(new_n738), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n732), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n789), .A2(new_n247), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n768), .B2(new_n829), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n758), .A2(new_n336), .B1(new_n779), .B2(new_n832), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n738), .B(new_n1002), .C1(G50), .C2(new_n830), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n772), .A2(new_n242), .B1(new_n751), .B2(new_n792), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n775), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(G58), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n758), .A2(new_n776), .B1(new_n779), .B2(new_n753), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n318), .B(new_n1008), .C1(G283), .C2(new_n830), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n772), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G107), .A2(new_n1010), .B1(new_n752), .B2(G294), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT46), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n775), .B2(new_n442), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n790), .A2(G97), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n782), .B2(new_n767), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n999), .B1(new_n1019), .B2(new_n746), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n960), .A2(new_n802), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n996), .A2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n670), .A2(new_n745), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n682), .A2(new_n734), .B1(G107), .B2(new_n207), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n682), .A2(KEYINPUT111), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n682), .A2(KEYINPUT111), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n263), .B1(new_n242), .B2(new_n247), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n382), .A2(new_n250), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(KEYINPUT50), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n739), .B1(new_n228), .B2(G45), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1025), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n747), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n732), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n827), .A2(G317), .B1(new_n830), .B2(G303), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n782), .B2(new_n751), .C1(new_n767), .C2(new_n757), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1010), .A2(G283), .B1(new_n1005), .B2(G294), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n790), .A2(G116), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n318), .B1(new_n780), .B2(new_n769), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n768), .A2(G159), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n758), .A2(new_n250), .B1(new_n783), .B2(new_n242), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n738), .B(new_n1051), .C1(G150), .C2(new_n780), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n772), .A2(new_n415), .B1(new_n751), .B2(new_n335), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n775), .A2(new_n247), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1052), .A3(new_n1016), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1036), .B1(new_n1057), .B2(new_n746), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n989), .A2(new_n731), .B1(new_n1024), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n990), .A2(new_n728), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n725), .A2(new_n989), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  NOR2_X1   g0862(.A1(new_n986), .A2(new_n990), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n683), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n986), .A2(new_n990), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n986), .A2(new_n730), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n747), .B1(new_n447), .B2(new_n207), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n238), .A2(new_n739), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1070), .A2(new_n733), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n767), .A2(new_n336), .B1(new_n792), .B2(new_n758), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1072), .B(new_n1073), .Z(new_n1074));
  NOR2_X1   g0874(.A1(new_n772), .A2(new_n247), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G50), .B2(new_n752), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n242), .B2(new_n775), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n318), .B1(new_n779), .B2(new_n828), .C1(new_n335), .C2(new_n783), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n837), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n767), .A2(new_n753), .B1(new_n782), .B2(new_n758), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n738), .B1(new_n779), .B2(new_n757), .C1(new_n773), .C2(new_n783), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G116), .A2(new_n1010), .B1(new_n752), .B2(G303), .ZN(new_n1083));
  INV_X1    g0883(.A(G283), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n775), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1082), .B(new_n1085), .C1(G107), .C2(new_n790), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1074), .A2(new_n1079), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1071), .B1(new_n749), .B2(new_n1087), .C1(new_n946), .C2(new_n802), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1066), .A2(new_n1067), .A3(new_n1088), .ZN(G390));
  OAI211_X1 g0889(.A(G330), .B(new_n932), .C1(new_n722), .C2(new_n723), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n694), .A2(new_n661), .A3(new_n817), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT115), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n891), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n713), .A2(new_n714), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n937), .B1(new_n1094), .B2(new_n721), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n817), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n889), .A2(KEYINPUT115), .A3(new_n890), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1090), .A2(new_n813), .A3(new_n1091), .A4(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n932), .A2(new_n1095), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n817), .C1(new_n722), .C2(new_n723), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n891), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n863), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n440), .A2(new_n1095), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n918), .A2(new_n639), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1091), .A2(new_n813), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT114), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n913), .B2(new_n914), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT102), .B1(new_n886), .B2(new_n667), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(KEYINPUT114), .A3(new_n912), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n926), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n667), .B(new_n816), .C1(new_n649), .C2(new_n651), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n813), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n891), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n909), .B1(new_n1123), .B2(new_n916), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n1124), .A3(new_n1090), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1093), .A2(new_n1097), .B1(new_n1091), .B2(new_n813), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1114), .B(new_n1116), .C1(new_n904), .C2(new_n906), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n907), .A2(new_n908), .B1(new_n1122), .B2(new_n915), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1100), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1109), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1105), .A2(new_n1125), .A3(new_n1130), .A4(new_n1108), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n728), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1125), .A2(new_n1130), .A3(new_n731), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n807), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n732), .B1(new_n382), .B2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n827), .A2(G116), .B1(new_n780), .B2(G294), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n447), .B2(new_n783), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1075), .B(new_n1139), .C1(G107), .C2(new_n752), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n738), .B1(new_n775), .B2(new_n589), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n768), .A2(G283), .B1(KEYINPUT117), .B2(new_n1141), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n819), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n318), .B1(new_n789), .B2(new_n250), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n768), .A2(G128), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n775), .A2(new_n336), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n783), .A2(new_n1150), .B1(new_n779), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G132), .B2(new_n827), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G159), .A2(new_n1010), .B1(new_n752), .B2(G137), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1147), .A2(new_n1149), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1137), .B1(new_n1156), .B2(new_n746), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n910), .B2(new_n744), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1134), .A2(new_n1159), .ZN(G378));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n892), .B1(new_n633), .B2(new_n660), .C1(new_n909), .C2(new_n915), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n344), .A2(new_n659), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n356), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n346), .B(new_n1163), .C1(new_n353), .C2(new_n355), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n934), .B2(G330), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n937), .B(new_n1173), .C1(new_n930), .C2(new_n933), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1162), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n932), .B(new_n922), .C1(new_n904), .C2(new_n906), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n929), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1178), .A2(KEYINPUT40), .B1(new_n1179), .B2(new_n931), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1173), .B1(new_n1180), .B2(new_n937), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n934), .A2(G330), .A3(new_n1174), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n917), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1161), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1107), .B(KEYINPUT119), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1133), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n683), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1177), .A2(new_n1183), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1189), .B2(KEYINPUT57), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n732), .B1(G50), .B2(new_n1136), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1174), .A2(new_n744), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n772), .A2(new_n336), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n827), .A2(G128), .B1(new_n830), .B2(G137), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n775), .B2(new_n1150), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(G132), .C2(new_n752), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1151), .B2(new_n767), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT118), .Z(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n790), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n790), .A2(G58), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n442), .B2(new_n767), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n738), .A2(new_n262), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G283), .B2(new_n780), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n514), .B2(new_n758), .C1(new_n415), .C2(new_n783), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1054), .B1(G68), .B2(new_n1010), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n447), .B2(new_n751), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1206), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT58), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1207), .B(new_n250), .C1(G33), .C2(G41), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1212), .A2(KEYINPUT58), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1204), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1191), .B(new_n1192), .C1(new_n1216), .C2(new_n746), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1188), .B2(new_n731), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1190), .A2(new_n1218), .ZN(G375));
  OAI211_X1 g1019(.A(new_n1107), .B(new_n1099), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1109), .A2(new_n993), .A3(new_n1220), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT120), .Z(new_n1222));
  NAND2_X1  g1022(.A1(new_n1105), .A2(new_n731), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n832), .A2(new_n758), .B1(new_n751), .B2(new_n1150), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n768), .B2(G132), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT123), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n318), .B1(new_n783), .B2(new_n336), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G128), .B2(new_n780), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1010), .A2(G50), .B1(new_n1005), .B2(G159), .ZN(new_n1229));
  AND4_X1   g1029(.A1(new_n1205), .A2(new_n1226), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n751), .A2(new_n442), .B1(new_n783), .B2(new_n514), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT121), .Z(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n773), .B2(new_n767), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n738), .B1(new_n779), .B2(new_n776), .C1(new_n447), .C2(new_n775), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n772), .A2(new_n415), .B1(new_n758), .B2(new_n1084), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT122), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1233), .A2(new_n1000), .A3(new_n1234), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n746), .B1(new_n1230), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n733), .B1(new_n242), .B2(new_n807), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n743), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1238), .B(new_n1239), .C1(new_n1110), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1223), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1222), .A2(new_n1243), .ZN(G381));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(G390), .A2(G384), .A3(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n975), .A2(new_n995), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  OR3_X1    g1049(.A1(new_n1249), .A2(G375), .A3(G381), .ZN(G407));
  INV_X1    g1050(.A(G375), .ZN(new_n1251));
  INV_X1    g1051(.A(G213), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(G343), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1248), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G407), .A2(G213), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT124), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT124), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(G407), .A2(new_n1257), .A3(G213), .A4(new_n1254), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(G409));
  XOR2_X1   g1059(.A(G393), .B(G396), .Z(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1247), .B2(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1260), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1262), .A2(new_n1263), .A3(G390), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1220), .B(KEYINPUT60), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n683), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1242), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(G384), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(G384), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G2897), .B(new_n1253), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1272), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(G384), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1253), .A2(G2897), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1189), .A2(new_n993), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1279), .B2(new_n1218), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n728), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1218), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT125), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1190), .A2(new_n1286), .A3(G378), .A4(new_n1218), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1280), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1278), .B1(new_n1288), .B2(new_n1253), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1253), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1267), .B(new_n1289), .C1(new_n1292), .C2(new_n1294), .ZN(new_n1295));
  XOR2_X1   g1095(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1296));
  NOR4_X1   g1096(.A1(new_n1288), .A2(new_n1253), .A3(new_n1291), .A4(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1266), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1253), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1280), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1278), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1303));
  INV_X1    g1103(.A(G390), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1262), .A2(new_n1263), .A3(G390), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1292), .A2(new_n1308), .ZN(new_n1309));
  NOR4_X1   g1109(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1291), .A4(new_n1253), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1302), .B(new_n1307), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1298), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(G378), .B2(new_n1251), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1290), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1314), .A2(new_n1290), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1307), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1314), .A2(new_n1290), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1266), .A2(new_n1315), .A3(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(G402));
endmodule


