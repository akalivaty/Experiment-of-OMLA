

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  XNOR2_X1 U322 ( .A(n344), .B(n343), .ZN(n347) );
  XNOR2_X1 U323 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U324 ( .A(n349), .B(n348), .ZN(n550) );
  XOR2_X1 U325 ( .A(KEYINPUT62), .B(n579), .Z(n290) );
  XOR2_X1 U326 ( .A(G211GAT), .B(G64GAT), .Z(n291) );
  XOR2_X1 U327 ( .A(KEYINPUT45), .B(n400), .Z(n292) );
  XNOR2_X1 U328 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n398) );
  XNOR2_X1 U329 ( .A(n399), .B(n398), .ZN(n403) );
  INV_X1 U330 ( .A(KEYINPUT11), .ZN(n341) );
  XNOR2_X1 U331 ( .A(n407), .B(n291), .ZN(n386) );
  XNOR2_X1 U332 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U333 ( .A(G99GAT), .B(G85GAT), .Z(n361) );
  NOR2_X1 U334 ( .A1(n565), .A2(n564), .ZN(n576) );
  NOR2_X1 U335 ( .A1(n523), .A2(n440), .ZN(n561) );
  XNOR2_X1 U336 ( .A(G183GAT), .B(KEYINPUT126), .ZN(n441) );
  XNOR2_X1 U337 ( .A(n442), .B(n441), .ZN(G1350GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n294) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(KEYINPUT80), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n312) );
  XOR2_X1 U341 ( .A(G190GAT), .B(G99GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U344 ( .A(G71GAT), .B(G120GAT), .Z(n298) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n310) );
  XOR2_X1 U348 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(G169GAT), .B(n303), .Z(n406) );
  XOR2_X1 U352 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n305) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n434) );
  XOR2_X1 U355 ( .A(n434), .B(G183GAT), .Z(n307) );
  NAND2_X1 U356 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n406), .B(n308), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X2 U360 ( .A(n312), .B(n311), .ZN(n523) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G106GAT), .Z(n336) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n314) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(G162GAT), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n422) );
  XOR2_X1 U365 ( .A(n336), .B(n422), .Z(n316) );
  NAND2_X1 U366 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U368 ( .A(G155GAT), .B(G204GAT), .Z(n318) );
  XNOR2_X1 U369 ( .A(G22GAT), .B(G148GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n320), .B(n319), .Z(n330) );
  XOR2_X1 U372 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n322) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(n323), .B(KEYINPUT85), .Z(n325) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G211GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n413) );
  XOR2_X1 U378 ( .A(G78GAT), .B(KEYINPUT22), .Z(n327) );
  XNOR2_X1 U379 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n413), .B(n328), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n454) );
  XOR2_X1 U383 ( .A(G43GAT), .B(KEYINPUT8), .Z(n332) );
  XNOR2_X1 U384 ( .A(KEYINPUT7), .B(KEYINPUT66), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n366) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n333), .B(KEYINPUT74), .ZN(n412) );
  XNOR2_X1 U388 ( .A(n366), .B(n412), .ZN(n349) );
  XOR2_X1 U389 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n335) );
  XNOR2_X1 U390 ( .A(G162GAT), .B(G92GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U392 ( .A(KEYINPUT72), .B(n361), .Z(n338) );
  XNOR2_X1 U393 ( .A(G218GAT), .B(n336), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(n340), .B(n339), .Z(n344) );
  NAND2_X1 U396 ( .A1(G232GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(G29GAT), .B(G134GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n345), .B(KEYINPUT73), .ZN(n433) );
  XNOR2_X1 U399 ( .A(n433), .B(KEYINPUT9), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n351) );
  XNOR2_X1 U402 ( .A(KEYINPUT69), .B(KEYINPUT32), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n354) );
  XNOR2_X1 U404 ( .A(G106GAT), .B(G57GAT), .ZN(n352) );
  XOR2_X1 U405 ( .A(G120GAT), .B(G148GAT), .Z(n428) );
  XNOR2_X1 U406 ( .A(n352), .B(n428), .ZN(n353) );
  XOR2_X1 U407 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U408 ( .A(G64GAT), .B(G92GAT), .Z(n356) );
  XNOR2_X1 U409 ( .A(G176GAT), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n410) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n357), .B(KEYINPUT13), .ZN(n392) );
  XNOR2_X1 U413 ( .A(n410), .B(n392), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U415 ( .A(n361), .B(n360), .Z(n363) );
  NAND2_X1 U416 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XOR2_X1 U417 ( .A(n363), .B(n362), .Z(n571) );
  XNOR2_X1 U418 ( .A(KEYINPUT41), .B(n571), .ZN(n540) );
  XOR2_X1 U419 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n365) );
  XNOR2_X1 U420 ( .A(G15GAT), .B(G22GAT), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n393) );
  XNOR2_X1 U422 ( .A(n366), .B(n393), .ZN(n379) );
  XOR2_X1 U423 ( .A(KEYINPUT29), .B(G8GAT), .Z(n368) );
  NAND2_X1 U424 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U426 ( .A(n369), .B(KEYINPUT30), .Z(n377) );
  XOR2_X1 U427 ( .A(G36GAT), .B(G50GAT), .Z(n371) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G29GAT), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U430 ( .A(G1GAT), .B(G141GAT), .Z(n373) );
  XNOR2_X1 U431 ( .A(G113GAT), .B(G197GAT), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n566) );
  INV_X1 U436 ( .A(n566), .ZN(n538) );
  NOR2_X1 U437 ( .A1(n540), .A2(n538), .ZN(n381) );
  XNOR2_X1 U438 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n396) );
  XOR2_X1 U440 ( .A(G57GAT), .B(G155GAT), .Z(n383) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(G127GAT), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n421) );
  XOR2_X1 U443 ( .A(KEYINPUT14), .B(n421), .Z(n385) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U446 ( .A(G8GAT), .B(G183GAT), .Z(n407) );
  XOR2_X1 U447 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n389) );
  XNOR2_X1 U448 ( .A(KEYINPUT76), .B(KEYINPUT12), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n391), .B(n390), .Z(n395) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n574) );
  XOR2_X1 U453 ( .A(KEYINPUT111), .B(n574), .Z(n528) );
  NOR2_X1 U454 ( .A1(n396), .A2(n528), .ZN(n397) );
  NAND2_X1 U455 ( .A1(n550), .A2(n397), .ZN(n399) );
  INV_X1 U456 ( .A(n574), .ZN(n545) );
  XNOR2_X1 U457 ( .A(n550), .B(KEYINPUT36), .ZN(n578) );
  NOR2_X1 U458 ( .A1(n545), .A2(n578), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n571), .A2(n292), .ZN(n401) );
  NAND2_X1 U460 ( .A1(n401), .A2(n538), .ZN(n402) );
  NAND2_X1 U461 ( .A1(n403), .A2(n402), .ZN(n405) );
  XOR2_X1 U462 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n519) );
  XOR2_X1 U464 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U465 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n506) );
  XNOR2_X1 U470 ( .A(KEYINPUT122), .B(n506), .ZN(n416) );
  NOR2_X1 U471 ( .A1(n519), .A2(n416), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n417), .B(KEYINPUT54), .ZN(n437) );
  XOR2_X1 U473 ( .A(KEYINPUT89), .B(KEYINPUT86), .Z(n419) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n420), .B(KEYINPUT1), .Z(n424) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT87), .Z(n426) );
  XNOR2_X1 U480 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U482 ( .A(n427), .B(KEYINPUT6), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(G85GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n459) );
  XNOR2_X1 U488 ( .A(KEYINPUT90), .B(n459), .ZN(n504) );
  NAND2_X1 U489 ( .A1(n437), .A2(n504), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n438), .B(KEYINPUT64), .ZN(n565) );
  NOR2_X1 U491 ( .A1(n454), .A2(n565), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n439), .B(KEYINPUT55), .ZN(n440) );
  NAND2_X1 U493 ( .A1(n561), .A2(n528), .ZN(n442) );
  NOR2_X1 U494 ( .A1(n571), .A2(n538), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n443), .B(KEYINPUT70), .ZN(n480) );
  XOR2_X1 U496 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n445) );
  NAND2_X1 U497 ( .A1(n574), .A2(n550), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n464) );
  XNOR2_X1 U499 ( .A(n506), .B(KEYINPUT27), .ZN(n450) );
  NOR2_X1 U500 ( .A1(n504), .A2(n450), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n446), .B(KEYINPUT91), .ZN(n518) );
  XOR2_X1 U502 ( .A(n454), .B(KEYINPUT65), .Z(n447) );
  XNOR2_X1 U503 ( .A(KEYINPUT28), .B(n447), .ZN(n474) );
  NOR2_X1 U504 ( .A1(n518), .A2(n474), .ZN(n448) );
  NAND2_X1 U505 ( .A1(n523), .A2(n448), .ZN(n462) );
  NAND2_X1 U506 ( .A1(n523), .A2(n454), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n449), .B(KEYINPUT26), .ZN(n564) );
  NOR2_X1 U508 ( .A1(n450), .A2(n564), .ZN(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT92), .B(n451), .Z(n457) );
  OR2_X1 U510 ( .A1(n523), .A2(n506), .ZN(n452) );
  XNOR2_X1 U511 ( .A(KEYINPUT93), .B(n452), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(KEYINPUT25), .B(n455), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U515 ( .A(KEYINPUT94), .B(n458), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n463), .B(KEYINPUT95), .ZN(n477) );
  NOR2_X1 U519 ( .A1(n464), .A2(n477), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT96), .ZN(n492) );
  NAND2_X1 U521 ( .A1(n480), .A2(n492), .ZN(n475) );
  NOR2_X1 U522 ( .A1(n504), .A2(n475), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U525 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U526 ( .A1(n506), .A2(n475), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(n469), .Z(n470) );
  XNOR2_X1 U528 ( .A(G8GAT), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U529 ( .A1(n523), .A2(n475), .ZN(n472) );
  XNOR2_X1 U530 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U532 ( .A(G15GAT), .B(n473), .Z(G1326GAT) );
  INV_X1 U533 ( .A(n474), .ZN(n521) );
  NOR2_X1 U534 ( .A1(n521), .A2(n475), .ZN(n476) );
  XOR2_X1 U535 ( .A(G22GAT), .B(n476), .Z(G1327GAT) );
  NOR2_X1 U536 ( .A1(n477), .A2(n578), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n545), .A2(n478), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT37), .ZN(n503) );
  NAND2_X1 U539 ( .A1(n480), .A2(n503), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT100), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT38), .B(n482), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n504), .A2(n490), .ZN(n485) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n483) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(n483), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  NOR2_X1 U546 ( .A1(n506), .A2(n490), .ZN(n486) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n486), .Z(G1329GAT) );
  NOR2_X1 U548 ( .A1(n523), .A2(n490), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U551 ( .A(G43GAT), .B(n489), .Z(G1330GAT) );
  NOR2_X1 U552 ( .A1(n521), .A2(n490), .ZN(n491) );
  XOR2_X1 U553 ( .A(G50GAT), .B(n491), .Z(G1331GAT) );
  NOR2_X1 U554 ( .A1(n566), .A2(n540), .ZN(n502) );
  NAND2_X1 U555 ( .A1(n502), .A2(n492), .ZN(n498) );
  NOR2_X1 U556 ( .A1(n504), .A2(n498), .ZN(n493) );
  XOR2_X1 U557 ( .A(G57GAT), .B(n493), .Z(n494) );
  XNOR2_X1 U558 ( .A(KEYINPUT42), .B(n494), .ZN(G1332GAT) );
  NOR2_X1 U559 ( .A1(n506), .A2(n498), .ZN(n496) );
  XNOR2_X1 U560 ( .A(G64GAT), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U561 ( .A(n496), .B(n495), .ZN(G1333GAT) );
  NOR2_X1 U562 ( .A1(n523), .A2(n498), .ZN(n497) );
  XOR2_X1 U563 ( .A(G71GAT), .B(n497), .Z(G1334GAT) );
  NOR2_X1 U564 ( .A1(n521), .A2(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U567 ( .A(G78GAT), .B(n501), .ZN(G1335GAT) );
  NAND2_X1 U568 ( .A1(n503), .A2(n502), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n504), .A2(n514), .ZN(n505) );
  XOR2_X1 U570 ( .A(G85GAT), .B(n505), .Z(G1336GAT) );
  NOR2_X1 U571 ( .A1(n506), .A2(n514), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G92GAT), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1337GAT) );
  NOR2_X1 U574 ( .A1(n523), .A2(n514), .ZN(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G99GAT), .B(n511), .ZN(G1338GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n513) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n516) );
  NOR2_X1 U581 ( .A1(n521), .A2(n514), .ZN(n515) );
  XOR2_X1 U582 ( .A(n516), .B(n515), .Z(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(n517), .ZN(G1339GAT) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(n520), .Z(n537) );
  NAND2_X1 U587 ( .A1(n521), .A2(n537), .ZN(n522) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n566), .A2(n532), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  INV_X1 U592 ( .A(n540), .ZN(n557) );
  NAND2_X1 U593 ( .A1(n532), .A2(n557), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n530) );
  NAND2_X1 U596 ( .A1(n532), .A2(n528), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n534) );
  INV_X1 U600 ( .A(n550), .ZN(n560) );
  NAND2_X1 U601 ( .A1(n532), .A2(n560), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n535), .ZN(G1343GAT) );
  INV_X1 U604 ( .A(n564), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n538), .A2(n549), .ZN(n539) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n539), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n549), .A2(n540), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n542) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n545), .A2(n549), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  XOR2_X1 U619 ( .A(G169GAT), .B(KEYINPUT123), .Z(n553) );
  NAND2_X1 U620 ( .A1(n561), .A2(n566), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n555) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(n556), .Z(n559) );
  NAND2_X1 U626 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT127), .Z(n568) );
  NAND2_X1 U632 ( .A1(n576), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n576), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U641 ( .A(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n290), .ZN(G1355GAT) );
endmodule

