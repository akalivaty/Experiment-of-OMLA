//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT87), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n202), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(G43gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n202), .B1(new_n208), .B2(KEYINPUT86), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n206), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n221), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n220), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT16), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n230), .A2(G1gat), .ZN(new_n234));
  OAI21_X1  g033(.A(G8gat), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n232), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n236), .B(new_n237), .C1(G1gat), .C2(new_n230), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n223), .A2(new_n229), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n238), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n241));
  INV_X1    g040(.A(new_n202), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n206), .A2(KEYINPUT87), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n208), .A2(new_n209), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n206), .A2(new_n225), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n208), .A2(KEYINPUT86), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n202), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n220), .B1(new_n249), .B2(new_n221), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n240), .B1(new_n251), .B2(KEYINPUT17), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(new_n246), .B2(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n239), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT18), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT18), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n223), .A2(new_n229), .A3(KEYINPUT17), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n235), .A2(new_n238), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n239), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n256), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n251), .A2(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n256), .B(KEYINPUT13), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G141gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G169gat), .B(G197gat), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT12), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n265), .A3(new_n269), .A4(new_n276), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT23), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n284), .A2(new_n286), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n291), .A2(KEYINPUT24), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT64), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT25), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT64), .B(new_n296), .C1(new_n290), .C2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(KEYINPUT65), .B2(KEYINPUT28), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT66), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n305), .A2(new_n282), .A3(new_n283), .A4(KEYINPUT66), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n289), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n302), .A2(new_n292), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n298), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(G120gat), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT68), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n314), .A2(new_n317), .A3(new_n320), .A4(new_n315), .ZN(new_n321));
  INV_X1    g120(.A(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G127gat), .ZN(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT1), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n329), .B2(KEYINPUT1), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n298), .A2(new_n331), .A3(new_n310), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G227gat), .ZN(new_n336));
  INV_X1    g135(.A(G233gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT34), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT32), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n336), .A2(new_n337), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n333), .A2(new_n341), .A3(new_n334), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n333), .A2(new_n344), .A3(new_n341), .A4(new_n334), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n340), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT33), .B1(new_n343), .B2(new_n345), .ZN(new_n347));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(KEYINPUT70), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(KEYINPUT70), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n353), .A2(KEYINPUT33), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n339), .B1(new_n351), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n338), .B(KEYINPUT34), .Z(new_n360));
  AND2_X1   g159(.A1(new_n343), .A2(new_n345), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n352), .B1(new_n361), .B2(new_n340), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n360), .B(new_n357), .C1(new_n362), .C2(new_n347), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT2), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n368), .B2(KEYINPUT2), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT73), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(G155gat), .B2(G162gat), .ZN(new_n374));
  INV_X1    g173(.A(G155gat), .ZN(new_n375));
  INV_X1    g174(.A(G162gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(G155gat), .A3(G162gat), .ZN(new_n380));
  AND4_X1   g179(.A1(new_n374), .A2(new_n377), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n376), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n368), .B1(new_n383), .B2(KEYINPUT2), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n367), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387));
  INV_X1    g186(.A(G211gat), .ZN(new_n388));
  INV_X1    g187(.A(G218gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n387), .B1(KEYINPUT22), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(KEYINPUT29), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n386), .B1(new_n394), .B2(KEYINPUT3), .ZN(new_n395));
  INV_X1    g194(.A(new_n393), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n372), .A2(new_n381), .B1(new_n367), .B2(new_n384), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G228gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n337), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n395), .B(new_n402), .C1(new_n396), .C2(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(G22gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(G22gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  NAND4_X1  g212(.A1(new_n408), .A2(new_n409), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n410), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n406), .B2(G22gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n413), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n415), .A2(new_n407), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n364), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n298), .A2(new_n310), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n298), .A2(new_n310), .B1(new_n425), .B2(new_n422), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n393), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n425), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n311), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n396), .A3(new_n423), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT71), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT71), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n434), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n427), .A2(new_n430), .ZN(new_n442));
  INV_X1    g241(.A(new_n433), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n397), .A2(new_n398), .B1(new_n328), .B2(new_n330), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(KEYINPUT5), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n328), .A2(new_n382), .A3(new_n385), .A4(new_n330), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n397), .A2(KEYINPUT76), .A3(new_n330), .A4(new_n328), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT4), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n458));
  INV_X1    g257(.A(new_n453), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n458), .B1(new_n457), .B2(new_n461), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n449), .B(new_n452), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT0), .ZN(new_n466));
  XNOR2_X1  g265(.A(G57gat), .B(G85gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n331), .A2(new_n386), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n456), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n471), .B2(new_n451), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT77), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n451), .B1(new_n447), .B2(new_n448), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT4), .B1(new_n455), .B2(new_n456), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n459), .A2(new_n460), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n464), .B(new_n468), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n472), .A2(new_n473), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n474), .A3(new_n479), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n468), .B1(new_n485), .B2(new_n464), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n464), .B1(new_n475), .B2(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(new_n468), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n488), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n446), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n486), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n489), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n482), .A3(new_n481), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT79), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n446), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n421), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n420), .A2(new_n500), .A3(new_n363), .A4(new_n359), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n499), .A2(new_n500), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n359), .A2(new_n363), .A3(KEYINPUT36), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT36), .B1(new_n359), .B2(new_n363), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n487), .A2(new_n490), .ZN(new_n506));
  INV_X1    g305(.A(new_n442), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n433), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT37), .B1(new_n430), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n507), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n434), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n442), .A2(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n510), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n419), .B1(new_n506), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n471), .A2(new_n451), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT82), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT39), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n521), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n449), .B1(new_n462), .B2(new_n463), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n451), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT39), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n527), .A3(new_n451), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n528), .A2(KEYINPUT81), .A3(new_n468), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT81), .B1(new_n528), .B2(new_n468), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT40), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n446), .A2(new_n486), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n526), .B(KEYINPUT40), .C1(new_n529), .C2(new_n530), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n505), .B1(new_n519), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n492), .A2(new_n419), .A3(new_n498), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n281), .B1(new_n502), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT90), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n542), .A2(KEYINPUT41), .ZN(new_n543));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT8), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  OR2_X1    g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G99gat), .B(G106gat), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G99gat), .B(G106gat), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n552), .C1(new_n557), .C2(new_n558), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n254), .A2(new_n259), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT8), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(G99gat), .B2(G106gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT91), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n556), .A3(new_n555), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n562), .B1(new_n571), .B2(new_n552), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n560), .B(new_n551), .C1(new_n569), .C2(new_n570), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n223), .A2(new_n229), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n542), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578));
  AND4_X1   g377(.A1(new_n565), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n574), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n542), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n580), .B2(new_n565), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n546), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(KEYINPUT93), .B(new_n546), .C1(new_n579), .C2(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n578), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n254), .A2(new_n259), .A3(new_n564), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n577), .B1(new_n251), .B2(new_n564), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n580), .A2(new_n565), .A3(new_n578), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n545), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT92), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n590), .A2(new_n594), .A3(new_n545), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n586), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G57gat), .B(G64gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT9), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n604), .B(new_n603), .C1(new_n599), .C2(new_n606), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  OAI21_X1  g413(.A(new_n260), .B1(new_n611), .B2(new_n610), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT88), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT89), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n620), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n616), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n563), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n610), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(new_n631), .C1(new_n572), .C2(new_n573), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n561), .B(new_n563), .C1(new_n629), .C2(new_n610), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n564), .A2(new_n635), .A3(new_n610), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n628), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n628), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G120gat), .B(G148gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT95), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n637), .B2(new_n639), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n627), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(KEYINPUT96), .A3(new_n644), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n540), .A2(new_n506), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g452(.A1(new_n540), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n446), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n237), .B2(new_n655), .ZN(new_n658));
  MUX2_X1   g457(.A(new_n657), .B(new_n658), .S(KEYINPUT42), .Z(G1325gat));
  OR2_X1    g458(.A1(new_n503), .A2(new_n504), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n359), .A2(new_n363), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(G15gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n654), .B2(new_n663), .ZN(G1326gat));
  NOR2_X1   g463(.A1(new_n654), .A2(new_n420), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT43), .B(G22gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NOR3_X1   g466(.A1(new_n650), .A2(new_n625), .A3(new_n281), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n536), .A2(new_n519), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n669), .A2(new_n538), .A3(new_n660), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n501), .A2(new_n491), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n662), .A2(new_n419), .ZN(new_n672));
  AOI211_X1 g471(.A(KEYINPUT79), .B(new_n445), .C1(new_n493), .C2(new_n495), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n497), .B1(new_n496), .B2(new_n446), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(KEYINPUT35), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n597), .B(new_n668), .C1(new_n670), .C2(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n677), .A2(G29gat), .A3(new_n496), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT45), .Z(new_n679));
  OAI211_X1 g478(.A(KEYINPUT44), .B(new_n597), .C1(new_n670), .C2(new_n676), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n668), .B(KEYINPUT97), .Z(new_n681));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n538), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n492), .A2(KEYINPUT98), .A3(new_n419), .A4(new_n498), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n537), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n598), .B1(new_n685), .B2(new_n502), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n680), .B(new_n681), .C1(new_n686), .C2(KEYINPUT44), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n496), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n679), .A2(new_n688), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n677), .A2(G36gat), .A3(new_n446), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n687), .B2(new_n446), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n687), .B2(new_n660), .ZN(new_n694));
  INV_X1    g493(.A(new_n650), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n662), .A2(G43gat), .A3(new_n598), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n540), .A2(new_n624), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT99), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT47), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  AOI211_X1 g500(.A(KEYINPUT99), .B(new_n701), .C1(new_n694), .C2(new_n697), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(G1330gat));
  OAI21_X1  g502(.A(G50gat), .B1(new_n687), .B2(new_n420), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n677), .A2(G50gat), .A3(new_n420), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1331gat));
  NAND2_X1  g507(.A1(new_n685), .A2(new_n502), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n626), .A2(new_n280), .A3(new_n695), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n506), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g513(.A1(new_n711), .A2(new_n446), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  AND2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n715), .B2(new_n716), .ZN(G1333gat));
  OAI21_X1  g518(.A(G71gat), .B1(new_n711), .B2(new_n660), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n364), .A2(new_n601), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n711), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT100), .B(KEYINPUT50), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1334gat));
  NOR2_X1   g523(.A1(new_n711), .A2(new_n420), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n602), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n625), .A2(new_n280), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT51), .B1(new_n686), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n727), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(KEYINPUT101), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n496), .A2(G85gat), .A3(new_n695), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT102), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n695), .A2(new_n280), .A3(new_n625), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n680), .B(new_n737), .C1(new_n686), .C2(KEYINPUT44), .ZN(new_n738));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738), .B2(new_n496), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(G1336gat));
  NOR3_X1   g539(.A1(new_n446), .A2(new_n695), .A3(G92gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n731), .A2(new_n733), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743));
  OAI21_X1  g542(.A(G92gat), .B1(new_n738), .B2(new_n446), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n730), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n741), .B1(new_n746), .B2(new_n728), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(G1337gat));
  NOR3_X1   g549(.A1(new_n662), .A2(G99gat), .A3(new_n695), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n731), .A2(new_n733), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G99gat), .B1(new_n738), .B2(new_n660), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1338gat));
  NOR3_X1   g553(.A1(new_n420), .A2(G106gat), .A3(new_n695), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n731), .A2(new_n733), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757));
  OAI21_X1  g556(.A(G106gat), .B1(new_n738), .B2(new_n420), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n746), .B2(new_n728), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n758), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1339gat));
  INV_X1    g562(.A(new_n643), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n637), .B2(KEYINPUT54), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n637), .A2(KEYINPUT54), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n634), .A2(new_n636), .A3(new_n628), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT103), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n632), .A2(new_n633), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n635), .ZN(new_n770));
  INV_X1    g569(.A(new_n636), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n638), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT103), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n772), .A2(new_n637), .A3(new_n773), .A4(KEYINPUT54), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n765), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n775), .A2(KEYINPUT55), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n645), .B1(new_n775), .B2(KEYINPUT55), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n280), .ZN(new_n778));
  INV_X1    g577(.A(new_n268), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n262), .A2(new_n266), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n256), .B1(new_n261), .B2(new_n262), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g582(.A(KEYINPUT104), .B(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n275), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n279), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT104), .B1(new_n255), .B2(new_n256), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n782), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(new_n780), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT105), .B1(new_n790), .B2(new_n275), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n650), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n597), .B1(new_n778), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n777), .A3(new_n597), .A4(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n624), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n651), .A2(new_n281), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n496), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n672), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n445), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n801), .A2(KEYINPUT107), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(KEYINPUT107), .ZN(new_n803));
  AOI211_X1 g602(.A(G113gat), .B(new_n281), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n419), .B1(new_n797), .B2(new_n798), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n496), .A2(new_n662), .A3(new_n445), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n281), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT106), .Z(new_n809));
  OR2_X1    g608(.A1(new_n804), .A2(new_n809), .ZN(G1340gat));
  NOR2_X1   g609(.A1(new_n695), .A2(G120gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n802), .B2(new_n803), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n814));
  INV_X1    g613(.A(new_n807), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n316), .B1(new_n815), .B2(new_n650), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n813), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1341gat));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n324), .A3(new_n625), .ZN(new_n820));
  OAI21_X1  g619(.A(G127gat), .B1(new_n807), .B2(new_n624), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT109), .ZN(G1342gat));
  NOR2_X1   g622(.A1(new_n598), .A2(new_n445), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n322), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n800), .A2(KEYINPUT110), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT110), .B1(new_n800), .B2(new_n825), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT111), .Z(new_n830));
  AOI21_X1  g629(.A(new_n322), .B1(new_n815), .B2(new_n597), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n828), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(KEYINPUT56), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1343gat));
  INV_X1    g633(.A(G141gat), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n496), .A2(new_n445), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n660), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n797), .A2(new_n798), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n838), .B2(new_n419), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n420), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n768), .A2(new_n774), .ZN(new_n842));
  INV_X1    g641(.A(new_n765), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n644), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n280), .B1(new_n775), .B2(KEYINPUT55), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n793), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n598), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n625), .B1(new_n848), .B2(new_n795), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n798), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT112), .B(new_n625), .C1(new_n848), .C2(new_n795), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n841), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n839), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT113), .B(new_n841), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n837), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n835), .B1(new_n857), .B2(new_n280), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n505), .A2(new_n420), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT114), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n281), .A2(G141gat), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n446), .A2(new_n860), .A3(new_n799), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT58), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  INV_X1    g663(.A(new_n799), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n660), .A2(new_n419), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n505), .A2(KEYINPUT114), .A3(new_n420), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT115), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n860), .A2(new_n871), .A3(new_n799), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n870), .A2(new_n872), .A3(new_n446), .A4(new_n861), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n864), .B1(new_n858), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n875), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n281), .B(new_n837), .C1(new_n855), .C2(new_n856), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n877), .B(KEYINPUT116), .C1(new_n835), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n876), .A3(new_n879), .ZN(G1344gat));
  NOR2_X1   g679(.A1(new_n695), .A2(G148gat), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n870), .A2(new_n872), .A3(new_n446), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT117), .Z(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n798), .B(KEYINPUT118), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n597), .B1(new_n775), .B2(KEYINPUT55), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n845), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n776), .A2(new_n777), .A3(KEYINPUT119), .A4(new_n597), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n792), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n848), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n625), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n848), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n840), .B1(new_n895), .B2(new_n420), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n838), .A2(new_n841), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n898), .A2(new_n660), .A3(new_n650), .A4(new_n836), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n884), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n884), .A2(G148gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n857), .B2(new_n650), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n883), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  AND2_X1   g702(.A1(new_n857), .A2(new_n625), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n870), .A2(new_n872), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n446), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n625), .A2(new_n375), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n904), .A2(new_n375), .B1(new_n906), .B2(new_n907), .ZN(G1346gat));
  NAND2_X1  g707(.A1(new_n857), .A2(new_n597), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n857), .A2(KEYINPUT121), .A3(new_n597), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(G162gat), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n905), .A2(new_n376), .A3(new_n824), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  NAND4_X1  g714(.A1(new_n805), .A2(new_n496), .A3(new_n445), .A4(new_n364), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(new_n282), .A3(new_n281), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n506), .B1(new_n797), .B2(new_n798), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n421), .A2(new_n446), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n280), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n282), .B2(new_n920), .ZN(G1348gat));
  OAI21_X1  g720(.A(G176gat), .B1(new_n916), .B2(new_n695), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n918), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n650), .A2(new_n283), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT122), .ZN(G1349gat));
  AND4_X1   g725(.A1(new_n299), .A2(new_n918), .A3(new_n625), .A4(new_n919), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n916), .B2(new_n624), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n916), .B2(new_n598), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(KEYINPUT61), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n597), .A2(new_n300), .ZN(new_n937));
  OAI221_X1 g736(.A(new_n936), .B1(KEYINPUT61), .B2(new_n935), .C1(new_n923), .C2(new_n937), .ZN(G1351gat));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n496), .A2(new_n445), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n505), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n896), .B2(new_n897), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n939), .B1(new_n944), .B2(new_n281), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(KEYINPUT126), .A3(new_n280), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(G197gat), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n918), .A2(new_n445), .A3(new_n859), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT125), .Z(new_n949));
  INV_X1    g748(.A(G197gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n950), .A3(new_n280), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n947), .A2(new_n951), .ZN(G1352gat));
  OAI21_X1  g751(.A(G204gat), .B1(new_n944), .B2(new_n695), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n948), .A2(G204gat), .A3(new_n695), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n388), .A3(new_n625), .ZN(new_n957));
  NAND2_X1  g756(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n388), .B1(new_n943), .B2(new_n625), .ZN(new_n959));
  NOR2_X1   g758(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AOI211_X1 g761(.A(new_n388), .B(new_n960), .C1(new_n943), .C2(new_n625), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  OAI21_X1  g763(.A(G218gat), .B1(new_n944), .B2(new_n598), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n389), .A3(new_n597), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1355gat));
endmodule


