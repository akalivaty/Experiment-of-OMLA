//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(new_n190), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT76), .B(G902), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G110), .B(G140), .ZN(new_n197));
  INV_X1    g011(.A(G227), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G953), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n197), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n209), .A2(new_n204), .A3(new_n203), .A4(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n216), .A3(G143), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n217), .A2(new_n218), .A3(G128), .A4(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n214), .A2(new_n216), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n224), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n221), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(KEYINPUT70), .B(new_n221), .C1(new_n223), .C2(new_n227), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT83), .B(G101), .Z(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G107), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n237));
  INV_X1    g051(.A(G107), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G104), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT82), .A2(G107), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT82), .A2(G107), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n239), .B1(new_n242), .B2(G104), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n233), .B(new_n237), .C1(new_n243), .C2(KEYINPUT3), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n234), .B1(new_n240), .B2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n236), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G101), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT82), .B(G107), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n235), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT84), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT10), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT0), .B(G128), .Z(new_n256));
  AOI21_X1  g070(.A(G143), .B1(new_n214), .B2(new_n216), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n225), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n217), .A2(KEYINPUT0), .A3(G128), .A4(new_n220), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT82), .A2(G107), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT82), .A2(G107), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(G104), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n239), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT3), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n262), .B(G101), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(G101), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n232), .A2(new_n255), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT86), .B(KEYINPUT10), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT1), .B1(new_n224), .B2(G146), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n217), .A2(new_n220), .B1(G128), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n221), .B1(new_n277), .B2(KEYINPUT85), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT64), .B(G146), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n219), .B1(new_n279), .B2(G143), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n276), .A2(G128), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n275), .B1(new_n284), .B2(new_n253), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n212), .B1(new_n273), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n252), .A2(new_n248), .ZN(new_n287));
  INV_X1    g101(.A(new_n233), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n267), .A2(new_n268), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(KEYINPUT10), .A3(new_n230), .A4(new_n231), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n270), .A2(new_n272), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n212), .A4(new_n285), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n200), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n200), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n277), .A2(KEYINPUT85), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n282), .B1(new_n280), .B2(new_n281), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n221), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n247), .B1(new_n246), .B2(G101), .ZN(new_n300));
  AOI211_X1 g114(.A(KEYINPUT84), .B(new_n251), .C1(new_n245), .C2(new_n236), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n302), .A3(new_n244), .ZN(new_n303));
  INV_X1    g117(.A(new_n228), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n287), .B2(new_n289), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT12), .B1(new_n306), .B2(new_n211), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT12), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n308), .B(new_n212), .C1(new_n303), .C2(new_n305), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n296), .B(new_n293), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n196), .B1(new_n295), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n194), .B1(new_n311), .B2(new_n193), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n293), .B1(new_n307), .B2(new_n309), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(KEYINPUT87), .B(new_n293), .C1(new_n307), .C2(new_n309), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n296), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n293), .A2(new_n296), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n291), .A2(new_n292), .ZN(new_n320));
  INV_X1    g134(.A(new_n285), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n211), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n318), .A2(new_n193), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n192), .B1(new_n313), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G116), .B(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G116), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n329), .A2(KEYINPUT5), .A3(G119), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT2), .B(G113), .Z(new_n333));
  AOI22_X1  g147(.A1(new_n328), .A2(new_n332), .B1(new_n333), .B2(new_n327), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n244), .A2(new_n248), .A3(new_n252), .A4(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n271), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n336));
  INV_X1    g150(.A(new_n327), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT2), .B(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n327), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT68), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT68), .B1(new_n339), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n269), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n335), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n345));
  XNOR2_X1  g159(.A(G110), .B(G122), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(new_n335), .C1(new_n336), .C2(new_n343), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT6), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n339), .A2(new_n340), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT68), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n272), .A3(new_n269), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n346), .B1(new_n356), .B2(new_n335), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT88), .B(new_n348), .C1(new_n350), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n344), .A2(new_n347), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT6), .A4(new_n349), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G953), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G224), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n260), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(new_n221), .C1(new_n223), .C2(new_n227), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT89), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(KEYINPUT89), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n368), .A2(KEYINPUT89), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n369), .A3(G224), .A4(new_n363), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n362), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n364), .A2(KEYINPUT7), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n368), .B(new_n379), .Z(new_n380));
  XNOR2_X1  g194(.A(new_n253), .B(new_n334), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n346), .B(KEYINPUT8), .Z(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(new_n349), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n383), .A2(new_n190), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n378), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n375), .B1(new_n358), .B2(new_n361), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n190), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(KEYINPUT90), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n366), .A2(KEYINPUT16), .A3(G140), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n396));
  AND2_X1   g210(.A1(KEYINPUT78), .A2(G140), .ZN(new_n397));
  NOR2_X1   g211(.A1(KEYINPUT78), .A2(G140), .ZN(new_n398));
  OAI21_X1  g212(.A(G125), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT79), .B1(new_n366), .B2(G140), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT79), .B(G125), .C1(new_n397), .C2(new_n398), .ZN(new_n402));
  AOI211_X1 g216(.A(KEYINPUT80), .B(new_n396), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT78), .A2(G140), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n366), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n400), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n402), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n404), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n395), .B1(new_n403), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n213), .ZN(new_n414));
  OAI211_X1 g228(.A(G146), .B(new_n395), .C1(new_n403), .C2(new_n412), .ZN(new_n415));
  INV_X1    g229(.A(G237), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n363), .A3(G214), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n224), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n416), .A2(new_n363), .A3(G143), .A4(G214), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n209), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT17), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n420), .B(new_n209), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n414), .A2(new_n415), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G113), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n234), .ZN(new_n428));
  NAND2_X1  g242(.A1(KEYINPUT18), .A2(G131), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n420), .B(new_n429), .Z(new_n430));
  XNOR2_X1  g244(.A(G125), .B(G140), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n279), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n411), .B2(new_n213), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n432), .C1(new_n411), .C2(new_n213), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n430), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n426), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n428), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n420), .B(new_n421), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n411), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n226), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n411), .A2(new_n404), .A3(KEYINPUT16), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n394), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n445), .B1(new_n449), .B2(G146), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n440), .B1(new_n450), .B2(new_n437), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n439), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(G475), .A2(G902), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT20), .ZN(new_n456));
  INV_X1    g270(.A(new_n453), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n439), .B2(new_n451), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT92), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT94), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n453), .B(KEYINPUT93), .Z(new_n462));
  AND4_X1   g276(.A1(new_n461), .A2(new_n452), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT20), .B1(new_n439), .B2(new_n451), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n461), .B1(new_n464), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n456), .B(new_n460), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(G116), .B(G122), .Z(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n249), .ZN(new_n468));
  XNOR2_X1  g282(.A(G128), .B(G143), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT13), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n224), .A2(G128), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n470), .B(G134), .C1(KEYINPUT13), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n202), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n469), .B(new_n202), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n329), .A2(KEYINPUT14), .A3(G122), .ZN(new_n476));
  OAI211_X1 g290(.A(G107), .B(new_n476), .C1(new_n467), .C2(KEYINPUT14), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n477), .C1(new_n249), .C2(new_n467), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G217), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n188), .A2(new_n480), .A3(G953), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT95), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n479), .B2(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G478), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n488), .A2(new_n195), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n488), .B2(new_n195), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G952), .ZN(new_n494));
  AOI211_X1 g308(.A(G953), .B(new_n494), .C1(G234), .C2(G237), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n363), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n439), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n428), .B1(new_n426), .B2(new_n438), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n190), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G475), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n466), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G214), .B1(G237), .B2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR4_X1   g320(.A1(new_n326), .A2(new_n393), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n355), .B1(new_n211), .B2(new_n261), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT66), .B1(new_n205), .B2(G134), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n202), .A3(G137), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n205), .A2(G134), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G131), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n210), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n513), .B2(G131), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n230), .A2(new_n518), .A3(new_n231), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT28), .B1(new_n508), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n211), .A2(new_n259), .A3(new_n258), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT69), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n211), .A2(new_n523), .A3(new_n259), .A4(new_n258), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n355), .ZN(new_n526));
  INV_X1    g340(.A(new_n355), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n519), .A2(new_n527), .A3(new_n522), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n520), .B1(new_n529), .B2(KEYINPUT28), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n416), .A2(new_n363), .A3(G210), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT27), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT29), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n196), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n539));
  INV_X1    g353(.A(new_n528), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n230), .A2(new_n518), .A3(new_n231), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n522), .A2(new_n524), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT30), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n513), .A2(G131), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT67), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n228), .A2(new_n545), .A3(new_n515), .A4(new_n210), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n546), .A2(new_n547), .A3(new_n521), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n540), .B1(new_n550), .B2(new_n355), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n534), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT29), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n521), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n355), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n528), .B2(new_n557), .ZN(new_n558));
  OR3_X1    g372(.A1(new_n558), .A2(new_n553), .A3(new_n520), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n538), .B(new_n539), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NOR2_X1   g379(.A1(G472), .A2(G902), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n548), .B1(new_n525), .B2(KEYINPUT30), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n534), .B(new_n528), .C1(new_n567), .C2(new_n527), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT71), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n553), .B1(new_n558), .B2(new_n520), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT74), .B(new_n553), .C1(new_n558), .C2(new_n520), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n576), .A3(KEYINPUT31), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT72), .B1(new_n568), .B2(KEYINPUT31), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n551), .A2(new_n580), .A3(new_n581), .A4(new_n534), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n565), .B(new_n566), .C1(new_n578), .C2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n582), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n586), .A2(new_n570), .A3(new_n577), .A4(new_n575), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n565), .B1(new_n587), .B2(new_n566), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n564), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n480), .B1(new_n195), .B2(G234), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT23), .ZN(new_n592));
  INV_X1    g406(.A(G119), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(G128), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n594), .B(new_n595), .C1(G119), .C2(new_n222), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G110), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT24), .B(G110), .Z(new_n598));
  XNOR2_X1  g412(.A(G119), .B(G128), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n447), .A2(new_n448), .ZN(new_n603));
  AOI21_X1  g417(.A(G146), .B1(new_n603), .B2(new_n395), .ZN(new_n604));
  INV_X1    g418(.A(new_n415), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n596), .A2(G110), .B1(new_n599), .B2(new_n598), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n432), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n415), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT22), .B(G137), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n363), .A2(G221), .A3(G234), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n610), .B(new_n611), .Z(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n601), .B1(new_n414), .B2(new_n415), .ZN(new_n615));
  INV_X1    g429(.A(new_n609), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n617), .A3(new_n195), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT25), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n591), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n590), .A2(G902), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n613), .A2(new_n617), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n621), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n507), .A2(new_n589), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n288), .ZN(G3));
  NAND2_X1  g441(.A1(new_n587), .A2(new_n195), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n566), .B1(new_n578), .B2(new_n583), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n284), .A2(new_n253), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n228), .B1(new_n302), .B2(new_n244), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n211), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n308), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n306), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT87), .B1(new_n636), .B2(new_n293), .ZN(new_n637));
  INV_X1    g451(.A(new_n317), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n200), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(G469), .A3(new_n323), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n191), .B1(new_n640), .B2(new_n312), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n625), .A2(new_n629), .A3(new_n630), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n466), .A2(new_n503), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n483), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n488), .A2(new_n644), .B1(new_n487), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(G478), .A3(new_n195), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n488), .A2(new_n195), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n489), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n506), .B1(new_n385), .B2(new_n389), .ZN(new_n652));
  INV_X1    g466(.A(new_n498), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  NAND2_X1  g472(.A1(new_n464), .A2(new_n453), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n456), .A2(new_n460), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n491), .A2(new_n492), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(G475), .B2(new_n502), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n653), .A2(new_n652), .A3(new_n660), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n238), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  INV_X1    g481(.A(new_n630), .ZN(new_n668));
  INV_X1    g482(.A(G472), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n587), .B2(new_n195), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n621), .A2(new_n622), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n606), .A2(new_n673), .A3(new_n609), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT97), .B1(new_n615), .B2(new_n616), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n614), .A2(KEYINPUT36), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n676), .B1(new_n674), .B2(new_n675), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n623), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT98), .ZN(new_n681));
  INV_X1    g495(.A(new_n676), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n673), .B1(new_n606), .B2(new_n609), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT97), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n677), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT98), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n623), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n672), .A2(new_n681), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n507), .A2(new_n671), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  XNOR2_X1  g506(.A(KEYINPUT99), .B(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n495), .B1(new_n496), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n662), .A2(new_n660), .A3(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n689), .A3(new_n652), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n589), .A2(new_n697), .A3(new_n641), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XNOR2_X1  g513(.A(new_n694), .B(KEYINPUT39), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n326), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n552), .A2(new_n534), .ZN(new_n704));
  INV_X1    g518(.A(new_n529), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(new_n553), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n669), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n585), .B2(new_n588), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT38), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n390), .A2(new_n710), .A3(new_n392), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n710), .B1(new_n390), .B2(new_n392), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n643), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n715), .A2(new_n689), .A3(new_n506), .A4(new_n661), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n703), .A2(new_n709), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n717), .B(KEYINPUT101), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  NAND2_X1  g533(.A1(new_n689), .A2(new_n652), .ZN(new_n720));
  INV_X1    g534(.A(new_n650), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n466), .B2(new_n503), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n695), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n589), .A3(new_n641), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  NAND2_X1  g540(.A1(new_n322), .A2(new_n293), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n727), .A2(new_n200), .B1(new_n319), .B2(new_n636), .ZN(new_n728));
  OAI21_X1  g542(.A(G469), .B1(new_n728), .B2(new_n196), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n311), .A2(new_n193), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n729), .A2(new_n730), .A3(new_n192), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n729), .A2(new_n730), .A3(new_n192), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT102), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n589), .A3(new_n625), .A4(new_n655), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n589), .A3(new_n625), .A4(new_n663), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NOR3_X1   g555(.A1(new_n720), .A2(new_n504), .A3(new_n734), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n589), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  OAI211_X1 g558(.A(new_n586), .B(new_n569), .C1(new_n534), .C2(new_n530), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n566), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n629), .A2(new_n625), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n643), .A2(new_n493), .A3(new_n652), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n661), .B1(new_n466), .B2(new_n503), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n652), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n733), .A2(new_n653), .A3(new_n735), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n747), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n747), .A2(new_n753), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  INV_X1    g574(.A(new_n723), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n628), .A2(G472), .B1(new_n566), .B2(new_n745), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n731), .A2(new_n652), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n689), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  NAND2_X1  g579(.A1(new_n393), .A2(new_n505), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n326), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n589), .A2(new_n767), .A3(new_n625), .A4(new_n761), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT42), .B1(new_n768), .B2(KEYINPUT105), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  AND3_X1   g587(.A1(new_n589), .A2(new_n767), .A3(new_n625), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n696), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  NAND3_X1  g590(.A1(new_n639), .A2(KEYINPUT45), .A3(new_n323), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n318), .B2(new_n324), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(G469), .ZN(new_n780));
  INV_X1    g594(.A(new_n194), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT106), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n781), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n730), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT106), .B1(new_n782), .B2(new_n783), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n192), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(new_n700), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT43), .B1(new_n643), .B2(new_n721), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT43), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n466), .A2(new_n792), .A3(new_n503), .A4(new_n650), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT107), .ZN(new_n795));
  INV_X1    g609(.A(new_n671), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n689), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n766), .B1(new_n798), .B2(KEYINPUT44), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n798), .A2(new_n800), .A3(KEYINPUT44), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT108), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n790), .B(new_n799), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n788), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT47), .B(new_n192), .C1(new_n786), .C2(new_n787), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n630), .A2(KEYINPUT32), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n810), .A2(new_n584), .B1(G472), .B2(new_n563), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n766), .A2(new_n723), .A3(new_n625), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n734), .A2(new_n505), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n712), .B2(new_n713), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n791), .A2(new_n495), .A3(new_n793), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n629), .A2(new_n625), .A3(new_n746), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n506), .B1(new_n390), .B2(new_n392), .ZN(new_n824));
  INV_X1    g638(.A(new_n495), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n734), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n824), .A2(new_n826), .A3(new_n625), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n707), .B1(new_n810), .B2(new_n584), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n643), .A2(new_n650), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT115), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n794), .A2(new_n825), .A3(new_n734), .A4(new_n766), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n689), .A3(new_n762), .ZN(new_n836));
  INV_X1    g650(.A(new_n819), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n731), .A2(new_n506), .ZN(new_n838));
  INV_X1    g652(.A(new_n713), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n838), .B1(new_n839), .B2(new_n711), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n747), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n823), .A2(new_n834), .A3(new_n836), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n819), .A2(new_n820), .A3(new_n766), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n729), .A2(new_n730), .A3(new_n191), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT113), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n807), .A2(new_n808), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n815), .B1(new_n848), .B2(KEYINPUT51), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n847), .A2(new_n844), .ZN(new_n851));
  OAI211_X1 g665(.A(KEYINPUT116), .B(new_n850), .C1(new_n851), .C2(new_n843), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n827), .A2(new_n828), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n494), .B(G953), .C1(new_n853), .C2(new_n722), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n589), .A2(new_n625), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n837), .A2(new_n747), .A3(new_n763), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n835), .A2(new_n855), .A3(new_n857), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n843), .A2(new_n850), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n807), .A2(new_n808), .A3(new_n845), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n844), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n862), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n849), .A2(new_n852), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n626), .A2(new_n690), .A3(new_n743), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n715), .A2(new_n493), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n651), .A2(KEYINPUT109), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT109), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n722), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n393), .A2(new_n506), .A3(new_n498), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n642), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n737), .A2(new_n740), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n759), .A2(new_n869), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n761), .A2(new_n762), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n660), .A2(new_n503), .A3(new_n661), .A4(new_n695), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n811), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n767), .A2(new_n689), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n774), .A2(new_n696), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n768), .A2(KEYINPUT105), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n886), .A3(new_n769), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n878), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n192), .B(new_n695), .C1(new_n313), .C2(new_n325), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n689), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n709), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n750), .A2(new_n751), .A3(new_n652), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n751), .B1(new_n750), .B2(new_n652), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n687), .B1(new_n686), .B2(new_n623), .ZN(new_n897));
  INV_X1    g711(.A(new_n623), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT98), .B(new_n898), .C1(new_n685), .C2(new_n677), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n641), .A2(new_n672), .A3(new_n900), .A4(new_n695), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n810), .A2(new_n584), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n708), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(KEYINPUT110), .A3(new_n753), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n725), .A2(new_n698), .A3(new_n764), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n905), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n888), .A2(new_n910), .A3(KEYINPUT53), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n876), .A2(new_n626), .A3(new_n690), .A4(new_n743), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n737), .A2(new_n740), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n772), .A3(new_n759), .A4(new_n883), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT111), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n908), .B2(new_n909), .ZN(new_n917));
  AND4_X1   g731(.A1(KEYINPUT110), .A2(new_n753), .A3(new_n709), .A4(new_n891), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT110), .B1(new_n903), .B2(new_n753), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n725), .A2(new_n698), .A3(new_n764), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT52), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n905), .A2(new_n907), .A3(new_n906), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(KEYINPUT111), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n915), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n868), .B(new_n911), .C1(new_n925), .C2(KEYINPUT53), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n888), .B2(new_n910), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n925), .B2(KEYINPUT53), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n867), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n494), .A2(new_n363), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n729), .A2(new_n730), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n506), .B(new_n191), .C1(new_n933), .C2(KEYINPUT49), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(new_n625), .C1(KEYINPUT49), .C2(new_n933), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n935), .A2(new_n714), .A3(new_n643), .A4(new_n721), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n828), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n932), .A2(KEYINPUT118), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G75));
  NOR2_X1   g756(.A1(new_n363), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n888), .A2(new_n910), .A3(KEYINPUT53), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n908), .A2(new_n909), .A3(new_n916), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT111), .B1(new_n922), .B2(new_n923), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n888), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT53), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n195), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT56), .B1(new_n951), .B2(new_n386), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n362), .B(new_n376), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT55), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n944), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  AOI211_X1 g770(.A(KEYINPUT56), .B(new_n954), .C1(new_n951), .C2(new_n386), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G51));
  OAI21_X1  g772(.A(new_n911), .B1(new_n925), .B2(KEYINPUT53), .ZN(new_n959));
  INV_X1    g773(.A(new_n868), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT119), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n926), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n959), .A2(KEYINPUT119), .A3(new_n960), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n194), .B(KEYINPUT57), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n728), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n780), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n959), .A2(new_n196), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT120), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n943), .B1(new_n968), .B2(new_n972), .ZN(G54));
  NAND3_X1  g787(.A1(new_n951), .A2(KEYINPUT58), .A3(G475), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n439), .A3(new_n451), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n951), .A2(KEYINPUT58), .A3(G475), .A4(new_n452), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n975), .A2(new_n976), .A3(new_n944), .ZN(G60));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT59), .Z(new_n979));
  NOR2_X1   g793(.A1(new_n948), .A2(new_n949), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT54), .B1(new_n980), .B2(new_n927), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n981), .B2(new_n926), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n944), .B1(new_n982), .B2(new_n646), .ZN(new_n983));
  INV_X1    g797(.A(new_n979), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n646), .A2(new_n963), .A3(new_n964), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n917), .A2(new_n924), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT53), .B1(new_n990), .B2(new_n888), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n686), .B(new_n989), .C1(new_n991), .C2(new_n945), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT121), .ZN(new_n993));
  INV_X1    g807(.A(new_n624), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n950), .B2(new_n988), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT121), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n959), .A2(new_n996), .A3(new_n686), .A4(new_n989), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n993), .A2(new_n944), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n992), .A2(KEYINPUT61), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n624), .B1(new_n959), .B2(new_n989), .ZN(new_n1002));
  NOR4_X1   g816(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT122), .A4(new_n943), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT122), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n992), .A2(KEYINPUT61), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n959), .A2(new_n989), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n943), .B1(new_n1006), .B2(new_n994), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1000), .B1(new_n1003), .B2(new_n1008), .ZN(G66));
  NAND2_X1  g823(.A1(new_n878), .A2(new_n363), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT123), .Z(new_n1011));
  INV_X1    g825(.A(G224), .ZN(new_n1012));
  OAI21_X1  g826(.A(G953), .B1(new_n497), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n358), .B(new_n361), .C1(G898), .C2(new_n363), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G69));
  INV_X1    g830(.A(G900), .ZN(new_n1017));
  OAI21_X1  g831(.A(G953), .B1(new_n198), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT125), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n550), .B(new_n444), .ZN(new_n1020));
  INV_X1    g834(.A(new_n874), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n700), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n774), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n813), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n804), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n907), .B(KEYINPUT124), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n718), .A2(KEYINPUT62), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n718), .A2(new_n1026), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT62), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1025), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1020), .B1(new_n1031), .B2(G953), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n855), .A2(new_n753), .ZN(new_n1034));
  OR3_X1    g848(.A1(new_n789), .A2(KEYINPUT126), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT126), .B1(new_n789), .B2(new_n1034), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n804), .A2(new_n1037), .A3(new_n1026), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n813), .A2(new_n772), .A3(new_n775), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n363), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1017), .A2(G953), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1020), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1019), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1019), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1044), .B(new_n1032), .C1(new_n1045), .C2(new_n1020), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1043), .A2(new_n1046), .ZN(G72));
  NOR2_X1   g861(.A1(new_n552), .A2(new_n534), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n1038), .A2(new_n878), .A3(new_n1039), .ZN(new_n1049));
  NAND2_X1  g863(.A1(G472), .A2(G902), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT63), .Z(new_n1051));
  INV_X1    g865(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1048), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g867(.A(new_n1048), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1054), .A2(new_n704), .A3(new_n1051), .ZN(new_n1055));
  OAI211_X1 g869(.A(new_n1053), .B(new_n944), .C1(new_n928), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1030), .A2(new_n1027), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1057), .A2(new_n804), .A3(new_n1024), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1051), .B1(new_n1058), .B2(new_n878), .ZN(new_n1059));
  OR2_X1    g873(.A1(new_n1059), .A2(KEYINPUT127), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n704), .B1(new_n1059), .B2(KEYINPUT127), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1056), .B1(new_n1060), .B2(new_n1061), .ZN(G57));
endmodule


