//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969;
  OAI21_X1  g000(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G71gat), .B(G78gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT95), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT21), .ZN(new_n209));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT90), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n215), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n218));
  OAI221_X1 g017(.A(KEYINPUT91), .B1(G1gat), .B2(new_n214), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(new_n208), .B2(KEYINPUT21), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n213), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G183gat), .B(G211gat), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n227), .B(new_n228), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n223), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n213), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G190gat), .B(G218gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  NOR2_X1   g036(.A1(G43gat), .A2(G50gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G43gat), .A2(G50gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT87), .B(G50gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n237), .B(new_n240), .C1(new_n242), .C2(G43gat), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n243), .A2(KEYINPUT88), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT14), .B(G29gat), .ZN(new_n245));
  INV_X1    g044(.A(G36gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT14), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n248), .A2(new_n246), .A3(G29gat), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n241), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n241), .B1(new_n243), .B2(KEYINPUT88), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n247), .A2(new_n249), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT17), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT17), .B1(new_n251), .B2(new_n254), .ZN(new_n260));
  NAND2_X1  g059(.A1(G85gat), .A2(G92gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n261), .B(new_n262), .Z(new_n263));
  NAND2_X1  g062(.A1(G99gat), .A2(G106gat), .ZN(new_n264));
  INV_X1    g063(.A(G85gat), .ZN(new_n265));
  INV_X1    g064(.A(G92gat), .ZN(new_n266));
  AOI22_X1  g065(.A1(KEYINPUT8), .A2(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G99gat), .B(G106gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n259), .A2(new_n260), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n270), .ZN(new_n273));
  NAND3_X1  g072(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n236), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT99), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT99), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n236), .C1(new_n272), .C2(new_n275), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT96), .ZN(new_n281));
  XNOR2_X1  g080(.A(G134gat), .B(G162gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n259), .A2(new_n260), .A3(new_n271), .ZN(new_n284));
  INV_X1    g083(.A(new_n236), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n285), .A3(new_n273), .A4(new_n274), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n277), .A2(new_n279), .A3(new_n283), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(new_n286), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n283), .B(KEYINPUT97), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n207), .ZN(new_n292));
  INV_X1    g091(.A(new_n208), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(new_n270), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n208), .A2(KEYINPUT10), .A3(new_n270), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G230gat), .A2(G233gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n294), .A2(new_n299), .ZN(new_n301));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G176gat), .B(G204gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n299), .B(KEYINPUT100), .Z(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(new_n296), .B2(new_n297), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n305), .B1(new_n309), .B2(new_n301), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n235), .A2(new_n291), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G148gat), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n319), .A2(new_n321), .B1(KEYINPUT2), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n322), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT74), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  OR2_X1    g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n322), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n323), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n320), .A2(G141gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n318), .A2(G148gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(KEYINPUT73), .A2(G155gat), .A3(G162gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n325), .B1(new_n336), .B2(new_n322), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G211gat), .A2(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT22), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G197gat), .A2(G204gat), .ZN(new_n343));
  AND2_X1   g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G211gat), .B(G218gat), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n342), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n351), .B2(new_n352), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n339), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n330), .A2(new_n338), .A3(new_n355), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n346), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n348), .B1(new_n342), .B2(new_n349), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n317), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n339), .A2(new_n351), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n317), .ZN(new_n368));
  INV_X1    g167(.A(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n360), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n358), .A2(KEYINPUT82), .A3(new_n359), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(G22gat), .B1(new_n365), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT74), .B1(new_n324), .B2(new_n325), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n328), .A2(new_n327), .A3(new_n322), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n334), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n322), .A2(new_n336), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n328), .A3(new_n335), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n323), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT3), .B1(new_n382), .B2(KEYINPUT81), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(new_n353), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n369), .B1(new_n358), .B2(new_n359), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n316), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n360), .A2(new_n370), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n363), .A3(new_n372), .ZN(new_n388));
  INV_X1    g187(.A(new_n368), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G22gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n393), .B(G50gat), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n374), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n374), .B2(new_n392), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n315), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n365), .A2(new_n373), .A3(G22gat), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n386), .B2(new_n390), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n374), .A2(new_n392), .A3(new_n395), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n314), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G127gat), .B(G134gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n407));
  INV_X1    g206(.A(G120gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G113gat), .ZN(new_n409));
  INV_X1    g208(.A(G113gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G120gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT1), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n407), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n409), .C2(new_n411), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n406), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT66), .B1(new_n417), .B2(KEYINPUT1), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(new_n419), .A3(new_n413), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n420), .A3(new_n405), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT23), .ZN(new_n424));
  NAND2_X1  g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT23), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(G169gat), .B2(G176gat), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(G183gat), .A2(G190gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n429), .A2(new_n430), .B1(new_n432), .B2(KEYINPUT65), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(KEYINPUT65), .B2(new_n432), .ZN(new_n438));
  AND4_X1   g237(.A1(KEYINPUT25), .A2(new_n424), .A3(new_n425), .A4(new_n427), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n423), .A2(KEYINPUT26), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n442), .B(new_n430), .C1(new_n444), .C2(new_n423), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT27), .B(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(G190gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT28), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT28), .B1(new_n447), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n422), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n416), .A2(new_n421), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n434), .A2(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n455));
  INV_X1    g254(.A(new_n451), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n445), .B1(new_n456), .B2(new_n449), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G227gat), .ZN(new_n460));
  INV_X1    g259(.A(G233gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT68), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n459), .A2(new_n462), .B1(new_n463), .B2(KEYINPUT34), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n462), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(KEYINPUT34), .ZN(new_n473));
  INV_X1    g272(.A(new_n462), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n453), .B2(new_n458), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(KEYINPUT33), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n472), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n472), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n464), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n476), .A2(new_n478), .ZN(new_n483));
  AOI221_X4 g282(.A(new_n477), .B1(KEYINPUT33), .B2(new_n471), .C1(new_n459), .C2(new_n462), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n463), .B(KEYINPUT34), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n464), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n472), .A2(new_n473), .A3(new_n479), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n404), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n455), .B2(new_n457), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n438), .A2(new_n439), .ZN(new_n492));
  INV_X1    g291(.A(new_n435), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n428), .B2(new_n433), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n452), .B(KEYINPUT70), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n495), .A3(new_n359), .ZN(new_n496));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n441), .A2(new_n452), .ZN(new_n502));
  INV_X1    g301(.A(new_n497), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n363), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n495), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n503), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n359), .A3(new_n497), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n363), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G8gat), .B(G36gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  NAND4_X1  g313(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT30), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n514), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n498), .A2(KEYINPUT71), .B1(new_n503), .B2(new_n502), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n369), .B1(new_n517), .B2(new_n501), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n510), .B(new_n516), .C1(new_n505), .C2(new_n363), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(KEYINPUT30), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n511), .A3(new_n514), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT72), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n520), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528));
  XOR2_X1   g327(.A(G1gat), .B(G29gat), .Z(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G85gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT5), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT76), .B1(new_n454), .B2(new_n339), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT76), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n381), .A2(new_n537), .A3(new_n421), .A4(new_n416), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n454), .A2(new_n339), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G225gat), .A2(G233gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n544), .A3(new_n538), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n367), .A2(KEYINPUT75), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n547), .B(KEYINPUT3), .C1(new_n377), .C2(new_n380), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(new_n454), .A3(new_n548), .A4(new_n358), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n422), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n545), .A2(new_n549), .A3(new_n541), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT4), .B1(new_n422), .B2(new_n381), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(KEYINPUT4), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n454), .A3(new_n358), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n547), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n535), .B(new_n541), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  AOI211_X1 g359(.A(new_n528), .B(new_n534), .C1(new_n552), .C2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n533), .B1(new_n555), .B2(new_n559), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT6), .B1(new_n562), .B2(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n552), .A2(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n533), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n489), .A2(new_n527), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n565), .B1(new_n563), .B2(KEYINPUT78), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT78), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n571), .B(KEYINPUT6), .C1(new_n562), .C2(new_n552), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n562), .A2(new_n552), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n528), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n563), .A2(KEYINPUT78), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n577), .A4(new_n565), .ZN(new_n578));
  INV_X1    g377(.A(new_n561), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n527), .A3(new_n489), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT35), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n581), .B2(KEYINPUT35), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n568), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n404), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n580), .B2(new_n527), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n482), .A2(KEYINPUT69), .A3(new_n488), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n482), .A2(KEYINPUT69), .A3(KEYINPUT36), .A4(new_n488), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT83), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT85), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n555), .A2(new_n549), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n542), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n597), .A2(new_n534), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT84), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n540), .A2(new_n542), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n544), .B1(new_n536), .B2(new_n538), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n556), .A2(new_n557), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n601), .A2(new_n602), .A3(new_n553), .ZN(new_n603));
  OAI211_X1 g402(.A(KEYINPUT39), .B(new_n600), .C1(new_n603), .C2(new_n541), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT40), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n597), .A3(new_n534), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT84), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n610), .A2(new_n565), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n594), .B1(new_n612), .B2(new_n527), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n565), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n608), .B2(new_n605), .ZN(new_n615));
  INV_X1    g414(.A(new_n520), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n522), .A2(new_n521), .A3(KEYINPUT30), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT72), .B1(new_n524), .B2(new_n525), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n619), .A3(KEYINPUT85), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n506), .A2(new_n511), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n516), .B1(new_n622), .B2(KEYINPUT37), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n363), .B1(new_n517), .B2(new_n501), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n508), .A2(new_n509), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT37), .B1(new_n626), .B2(new_n369), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n624), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n566), .B(new_n524), .C1(new_n623), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n516), .A2(KEYINPUT37), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n519), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n622), .A2(KEYINPUT37), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n586), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n593), .B1(new_n621), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n590), .A2(new_n591), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n580), .A2(new_n527), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(new_n586), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT83), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n585), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n259), .A2(new_n221), .A3(new_n260), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n257), .A2(new_n222), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT92), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT18), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n641), .A2(KEYINPUT18), .A3(new_n642), .A4(new_n643), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n257), .B(new_n222), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n642), .B(KEYINPUT13), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G113gat), .B(G141gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G197gat), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT11), .B(G169gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT12), .Z(new_n659));
  NOR2_X1   g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n653), .A3(new_n650), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n659), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n640), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n313), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n580), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT101), .B(G1gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  INV_X1    g472(.A(new_n669), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT16), .B(G8gat), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n674), .A2(new_n527), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n220), .B1(new_n669), .B2(new_n619), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT42), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(KEYINPUT42), .B2(new_n676), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n674), .B2(new_n636), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n482), .A2(new_n488), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n674), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n669), .A2(new_n404), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NOR2_X1   g485(.A1(new_n235), .A2(new_n311), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n287), .A2(new_n290), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n693), .A2(G29gat), .A3(new_n580), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n634), .B1(new_n613), .B2(new_n620), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n638), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n698), .B(new_n568), .C1(new_n583), .C2(new_n584), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT86), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT35), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n698), .B1(new_n704), .B2(new_n568), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n688), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n291), .A2(new_n707), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n706), .A2(new_n707), .B1(new_n640), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n665), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n235), .A3(new_n311), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n580), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n713), .ZN(G1328gat));
  NAND2_X1  g513(.A1(new_n619), .A2(new_n246), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n693), .A2(new_n715), .B1(KEYINPUT103), .B2(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n712), .B2(new_n527), .ZN(new_n719));
  OAI211_X1 g518(.A(KEYINPUT103), .B(KEYINPUT46), .C1(new_n693), .C2(new_n715), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT104), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n718), .A2(new_n723), .A3(new_n719), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1329gat));
  OAI21_X1  g524(.A(G43gat), .B1(new_n712), .B2(new_n636), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n689), .B1(new_n667), .B2(new_n668), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n681), .A2(G43gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n726), .B(new_n729), .C1(KEYINPUT105), .C2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1330gat));
  NOR2_X1   g531(.A1(new_n586), .A2(new_n242), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n693), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n709), .A2(new_n404), .A3(new_n711), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n242), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n738), .ZN(new_n741));
  OAI221_X1 g540(.A(KEYINPUT48), .B1(new_n735), .B2(new_n736), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n735), .A2(new_n736), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n737), .A2(new_n242), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(KEYINPUT48), .B2(new_n745), .ZN(G1331gat));
  NAND4_X1  g545(.A1(new_n710), .A2(new_n235), .A3(new_n291), .A4(new_n311), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n638), .A2(new_n696), .ZN(new_n748));
  INV_X1    g547(.A(new_n568), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n702), .B2(new_n703), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(new_n698), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n585), .A2(KEYINPUT102), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n670), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT108), .B(G57gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1332gat));
  XNOR2_X1  g555(.A(new_n619), .B(KEYINPUT109), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT110), .ZN(G1333gat));
  NAND2_X1  g562(.A1(new_n753), .A2(new_n592), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n681), .A2(G71gat), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n764), .A2(G71gat), .B1(new_n753), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n753), .A2(new_n404), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT111), .B(G78gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n235), .A2(new_n665), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n709), .A2(new_n311), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n580), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(new_n688), .C1(new_n700), .C2(new_n705), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n771), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n752), .A2(new_n699), .A3(new_n697), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n774), .B1(new_n777), .B2(new_n688), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(KEYINPUT113), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n776), .B2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n706), .A2(KEYINPUT112), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(KEYINPUT51), .A3(new_n771), .A4(new_n775), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n670), .A2(new_n265), .A3(new_n311), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n773), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(G92gat), .B1(new_n772), .B2(new_n757), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n757), .A2(G92gat), .A3(new_n312), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n790), .B(new_n791), .C1(new_n787), .C2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n771), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n291), .B1(new_n751), .B2(new_n752), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n774), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n797), .B2(new_n783), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n792), .B1(new_n798), .B2(new_n780), .ZN(new_n799));
  OAI21_X1  g598(.A(G92gat), .B1(new_n772), .B2(new_n527), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n801), .B2(KEYINPUT52), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n793), .B1(new_n782), .B2(new_n784), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n771), .A2(new_n311), .ZN(new_n804));
  AOI221_X4 g603(.A(new_n804), .B1(new_n640), .B2(new_n708), .C1(new_n706), .C2(new_n707), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n266), .B1(new_n805), .B2(new_n619), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n803), .C2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n794), .B1(new_n802), .B2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n772), .B2(new_n636), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n681), .A2(G99gat), .A3(new_n312), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n787), .B2(new_n811), .ZN(G1338gat));
  INV_X1    g611(.A(G106gat), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n805), .B2(new_n404), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n312), .A2(new_n586), .A3(G106gat), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n787), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n798), .B2(new_n780), .ZN(new_n819));
  OAI21_X1  g618(.A(G106gat), .B1(new_n772), .B2(new_n586), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT115), .B1(new_n821), .B2(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n817), .B1(new_n782), .B2(new_n784), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n823), .C2(new_n814), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n818), .B1(new_n822), .B2(new_n825), .ZN(G1339gat));
  NOR2_X1   g625(.A1(new_n313), .A2(new_n665), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n642), .B1(new_n641), .B2(new_n643), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(new_n651), .B2(new_n652), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n658), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n291), .A2(new_n661), .A3(new_n311), .A4(new_n832), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n287), .A2(new_n290), .B1(new_n649), .B2(new_n660), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n834), .A2(new_n832), .B1(new_n665), .B2(new_n291), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n304), .B1(new_n309), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n298), .B2(new_n299), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n296), .A2(new_n308), .A3(new_n297), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT116), .B1(new_n839), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n843), .A2(new_n844), .B1(new_n300), .B2(new_n306), .ZN(new_n845));
  OAI211_X1 g644(.A(KEYINPUT55), .B(new_n837), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n833), .B1(new_n835), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n235), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n827), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n404), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n580), .A2(new_n681), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n758), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n710), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n665), .A2(new_n410), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT120), .Z(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n857), .B2(new_n860), .ZN(G1340gat));
  NOR2_X1   g660(.A1(new_n857), .A2(new_n312), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(new_n408), .ZN(G1341gat));
  NOR2_X1   g662(.A1(new_n857), .A2(new_n852), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(new_n212), .ZN(G1342gat));
  NAND2_X1  g664(.A1(new_n688), .A2(new_n527), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n855), .A3(G134gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT56), .Z(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n857), .B2(new_n291), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  OAI21_X1  g670(.A(KEYINPUT57), .B1(new_n853), .B2(new_n586), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n636), .A2(new_n670), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n758), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n846), .B(new_n847), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n688), .A2(new_n832), .A3(new_n661), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n688), .B1(new_n664), .B2(new_n661), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n876), .B(new_n845), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n235), .B1(new_n879), .B2(new_n833), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n875), .B(new_n404), .C1(new_n880), .C2(new_n827), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT121), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n872), .A2(new_n881), .A3(new_n884), .A4(new_n874), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n665), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n853), .A2(new_n586), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n874), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n710), .A2(G141gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT58), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n886), .A2(G141gat), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n882), .B2(new_n710), .ZN(new_n898));
  XOR2_X1   g697(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n898), .A2(KEYINPUT124), .A3(new_n891), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n894), .A2(new_n897), .A3(new_n904), .ZN(G1344gat));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n320), .A3(new_n311), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n883), .A2(new_n311), .A3(new_n885), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .A3(new_n320), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n872), .A2(new_n881), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n874), .A2(KEYINPUT125), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n874), .A2(KEYINPUT125), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n311), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G148gat), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n906), .B1(new_n908), .B2(new_n914), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n889), .A2(new_n226), .A3(new_n235), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n883), .A2(new_n235), .A3(new_n885), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n226), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n883), .A2(new_n688), .A3(new_n885), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G162gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n873), .A2(G162gat), .A3(new_n866), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n888), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n853), .A2(new_n670), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n619), .A3(new_n489), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n710), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n924), .A2(new_n489), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n758), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n928), .A2(G169gat), .A3(new_n710), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(G1348gat));
  OAI21_X1  g731(.A(G176gat), .B1(new_n925), .B2(new_n312), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n312), .A2(G176gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n928), .B2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n925), .B2(new_n852), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n235), .A2(new_n447), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n925), .B2(new_n291), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n688), .A2(new_n448), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n944), .A2(new_n945), .B1(new_n928), .B2(new_n946), .ZN(G1351gat));
  INV_X1    g746(.A(new_n909), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n592), .A2(new_n670), .A3(new_n527), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n950), .A2(new_n951), .A3(new_n710), .ZN(new_n952));
  AND4_X1   g751(.A1(new_n404), .A2(new_n924), .A3(new_n636), .A4(new_n758), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n665), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n952), .A2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n956), .A3(new_n311), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n950), .B2(new_n312), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1353gat));
  INV_X1    g759(.A(G211gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(new_n961), .A3(new_n235), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n948), .A2(new_n235), .A3(new_n949), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n950), .B2(new_n291), .ZN(new_n967));
  INV_X1    g766(.A(G218gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n968), .A3(new_n688), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1355gat));
endmodule


