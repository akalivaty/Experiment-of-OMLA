//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G134), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT11), .A2(G134), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT67), .B1(new_n198), .B2(new_n191), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT11), .A2(G134), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n200), .A2(new_n201), .A3(G137), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n195), .B(new_n197), .C1(new_n199), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(KEYINPUT67), .A3(new_n191), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n201), .B1(new_n200), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT68), .B(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(new_n195), .A4(new_n197), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT64), .A2(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(G143), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n212), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n215), .A2(new_n218), .A3(G128), .A4(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n214), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n225), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n221), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT10), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT87), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT87), .A2(G104), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT3), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n231), .A3(G104), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT88), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n236), .A2(new_n231), .A3(KEYINPUT88), .A4(G104), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  OR3_X1    g056(.A1(new_n232), .A2(new_n233), .A3(new_n231), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n235), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n234), .B1(G104), .B2(new_n231), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n230), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n228), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT64), .A2(G146), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT64), .A2(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n219), .B1(new_n253), .B2(G143), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT0), .A4(G128), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n215), .A2(KEYINPUT0), .A3(G128), .A4(new_n220), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n250), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n235), .A2(new_n243), .ZN(new_n261));
  INV_X1    g075(.A(new_n241), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n260), .B(G101), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n244), .A2(KEYINPUT4), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n232), .A2(new_n233), .A3(new_n231), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(KEYINPUT3), .B2(new_n234), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n242), .B1(new_n267), .B2(new_n241), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n248), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n226), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n222), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n221), .B1(new_n254), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n244), .A3(new_n246), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT89), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n274), .A2(new_n244), .A3(new_n277), .A4(new_n246), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n210), .B1(new_n271), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n259), .A2(new_n263), .ZN(new_n283));
  OAI22_X1  g097(.A1(new_n283), .A2(new_n269), .B1(new_n247), .B2(new_n230), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT10), .B1(new_n276), .B2(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n204), .A2(new_n209), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n190), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n281), .A3(new_n210), .ZN(new_n289));
  INV_X1    g103(.A(new_n190), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n229), .B1(new_n244), .B2(new_n246), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n279), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT12), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n276), .B2(new_n278), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT12), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(new_n210), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n289), .B(new_n290), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n286), .B1(new_n284), .B2(new_n285), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n289), .A2(new_n303), .A3(new_n290), .ZN(new_n304));
  INV_X1    g118(.A(new_n297), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n296), .B1(new_n295), .B2(new_n210), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n287), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n190), .B(KEYINPUT86), .ZN(new_n308));
  OAI211_X1 g122(.A(G469), .B(new_n304), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G469), .A2(G902), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n302), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  OAI21_X1  g126(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT90), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G119), .ZN(new_n320));
  INV_X1    g134(.A(G119), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT71), .A3(G116), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(G119), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT2), .B(G113), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT5), .A4(new_n323), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n319), .A2(KEYINPUT5), .A3(G119), .ZN(new_n329));
  INV_X1    g143(.A(G113), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n325), .A2(new_n327), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n244), .A3(new_n246), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n324), .B(new_n326), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n263), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n269), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n337), .B(new_n333), .C1(new_n269), .C2(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n221), .C1(new_n224), .C2(new_n228), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n250), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n348), .B2(G125), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G224), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n343), .B1(new_n259), .B2(new_n342), .ZN(new_n353));
  INV_X1    g167(.A(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n336), .A2(new_n357), .A3(new_n338), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n341), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT91), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n337), .B(KEYINPUT8), .ZN(new_n364));
  INV_X1    g178(.A(new_n333), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n332), .B1(new_n244), .B2(new_n246), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n355), .A2(new_n340), .A3(new_n363), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n351), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n301), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n359), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n361), .ZN(new_n373));
  AND4_X1   g187(.A1(new_n355), .A2(new_n340), .A3(new_n363), .A4(new_n367), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n374), .B2(new_n369), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n341), .A2(new_n356), .A3(new_n358), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n317), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n361), .B1(new_n359), .B2(new_n371), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n373), .A3(new_n376), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT92), .A3(new_n317), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n314), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n386));
  INV_X1    g200(.A(new_n208), .ZN(new_n387));
  OR2_X1    g201(.A1(KEYINPUT72), .A2(G237), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT72), .A2(G237), .ZN(new_n389));
  AOI21_X1  g203(.A(G953), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G143), .B1(new_n390), .B2(G214), .ZN(new_n391));
  AND2_X1   g205(.A1(KEYINPUT72), .A2(G237), .ZN(new_n392));
  NOR2_X1   g206(.A1(KEYINPUT72), .A2(G237), .ZN(new_n393));
  OAI211_X1 g207(.A(G214), .B(new_n350), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n225), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n387), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(G143), .A3(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n225), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n208), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n342), .B2(G140), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT76), .B(G140), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n342), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT76), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G140), .ZN(new_n406));
  INV_X1    g220(.A(G140), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT76), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n401), .B(G125), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(KEYINPUT19), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n342), .A2(G140), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g227(.A1(KEYINPUT94), .A2(KEYINPUT19), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT94), .A2(KEYINPUT19), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n253), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n400), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT78), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n404), .A2(new_n409), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT16), .ZN(new_n422));
  AOI211_X1 g236(.A(KEYINPUT78), .B(new_n422), .C1(new_n404), .C2(new_n409), .ZN(new_n423));
  OAI21_X1  g237(.A(G146), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n394), .B(G143), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT18), .B(G131), .C1(new_n391), .C2(new_n395), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n404), .A2(G146), .A3(new_n409), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n413), .A2(new_n253), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(KEYINPUT93), .A3(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n418), .A2(new_n424), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT95), .B(G104), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n386), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n430), .A2(KEYINPUT93), .A3(new_n431), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT93), .B1(new_n430), .B2(new_n431), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n427), .B(new_n428), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n420), .A2(KEYINPUT16), .ZN(new_n446));
  INV_X1    g260(.A(new_n419), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n412), .A2(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n407), .A2(KEYINPUT76), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n405), .A2(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n450), .B1(new_n453), .B2(G125), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n403), .A2(KEYINPUT77), .A3(new_n342), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n449), .B(KEYINPUT16), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n212), .B1(new_n448), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n400), .A2(new_n417), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n445), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT96), .A3(new_n440), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n442), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n422), .B1(new_n404), .B2(new_n409), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n456), .B(new_n212), .C1(new_n462), .C2(new_n419), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n424), .A2(KEYINPUT79), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(G146), .C1(new_n421), .C2(new_n423), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n396), .A2(new_n468), .A3(new_n399), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n396), .A2(KEYINPUT97), .A3(new_n468), .A4(new_n399), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n396), .A2(new_n468), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n441), .A3(new_n445), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n461), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g291(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT98), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n424), .A2(new_n400), .A3(new_n417), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n386), .B(new_n441), .C1(new_n481), .C2(new_n445), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT96), .B1(new_n459), .B2(new_n440), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n445), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n440), .B(new_n485), .C1(new_n467), .C2(new_n474), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n480), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n461), .A2(KEYINPUT98), .A3(new_n476), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n479), .B1(new_n490), .B2(KEYINPUT20), .ZN(new_n491));
  INV_X1    g305(.A(G475), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n441), .B1(new_n475), .B2(new_n445), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n494), .B2(new_n301), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n225), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n222), .A2(G143), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G134), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(G116), .B(G122), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n231), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n319), .A2(KEYINPUT14), .A3(G122), .ZN(new_n503));
  INV_X1    g317(.A(new_n501), .ZN(new_n504));
  OAI211_X1 g318(.A(G107), .B(new_n503), .C1(new_n504), .C2(KEYINPUT14), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n496), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n507), .A2(KEYINPUT13), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n497), .B1(new_n507), .B2(KEYINPUT13), .ZN(new_n509));
  OAI21_X1  g323(.A(G134), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n498), .A2(new_n499), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n501), .B(new_n231), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G217), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n312), .A2(new_n515), .A3(G953), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n514), .B(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n518), .A2(new_n301), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G478), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n520), .A3(new_n301), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n523), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(G234), .A2(G237), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n528), .A2(G952), .A3(new_n350), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT100), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n528), .A2(G902), .A3(G953), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n524), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n491), .A2(new_n495), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n385), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n390), .A2(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT27), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G101), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n334), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n256), .A2(new_n258), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n286), .A2(new_n546), .A3(new_n345), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n191), .A2(KEYINPUT69), .A3(G134), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n197), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT69), .B1(new_n191), .B2(G134), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n229), .A2(new_n209), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n545), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n209), .A2(new_n551), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n259), .A2(new_n286), .B1(new_n555), .B2(new_n229), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n545), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n544), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n552), .B1(new_n348), .B2(new_n210), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(new_n334), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n543), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n544), .B1(new_n556), .B2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n562), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n556), .A2(new_n544), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT28), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n568), .A3(new_n542), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n561), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT74), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n561), .A2(new_n569), .A3(new_n573), .A4(new_n570), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT29), .A4(new_n542), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n301), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n547), .A2(new_n545), .A3(new_n552), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n334), .B1(new_n580), .B2(new_n553), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n556), .A2(new_n544), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n542), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT31), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n334), .B1(new_n559), .B2(new_n564), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT28), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n559), .A2(new_n334), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n562), .B1(new_n588), .B2(new_n582), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n543), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(new_n591), .A3(new_n542), .A4(new_n582), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n584), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT32), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT32), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n595), .A2(KEYINPUT75), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n579), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(G119), .B(G128), .Z(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT24), .B(G110), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n321), .B2(G128), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n606), .B(new_n607), .C1(G119), .C2(new_n222), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(G110), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n464), .A2(new_n466), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n602), .A2(new_n603), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n608), .B2(G110), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT80), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n431), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n613), .B2(new_n612), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n424), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT82), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT22), .B(G137), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(G902), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT81), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n610), .A2(new_n624), .A3(new_n616), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n610), .B2(new_n616), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n620), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT83), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n610), .A2(new_n616), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT81), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n610), .A2(new_n624), .A3(new_n616), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(KEYINPUT83), .A3(new_n632), .A4(new_n628), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n623), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT25), .ZN(new_n636));
  INV_X1    g450(.A(new_n623), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n631), .A2(new_n632), .A3(new_n628), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT83), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n637), .B1(new_n640), .B2(new_n633), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT25), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n515), .B1(G234), .B2(new_n301), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n636), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n644), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n623), .B(new_n646), .C1(new_n629), .C2(new_n634), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(KEYINPUT84), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT84), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n641), .B2(new_n646), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n601), .A2(KEYINPUT85), .A3(new_n645), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n647), .A2(KEYINPUT84), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n641), .A2(new_n649), .A3(new_n646), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n644), .B1(new_n641), .B2(new_n642), .ZN(new_n656));
  AOI211_X1 g470(.A(KEYINPUT25), .B(new_n637), .C1(new_n640), .C2(new_n633), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n576), .B1(new_n571), .B2(KEYINPUT74), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n574), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n593), .A2(new_n594), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT32), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT75), .A3(new_n595), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n596), .A2(new_n598), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n653), .B1(new_n658), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n538), .B1(new_n652), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n242), .ZN(G3));
  INV_X1    g484(.A(new_n658), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n593), .A2(new_n301), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G472), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n313), .A2(new_n311), .A3(new_n673), .A4(new_n662), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n490), .A2(KEYINPUT20), .ZN(new_n676));
  INV_X1    g490(.A(new_n479), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n495), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT33), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(KEYINPUT102), .ZN(new_n683));
  MUX2_X1   g497(.A(new_n681), .B(new_n683), .S(new_n518), .Z(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(G478), .A3(new_n301), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(G478), .B2(new_n519), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n355), .A2(new_n367), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n369), .A3(new_n340), .A4(new_n363), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n376), .A2(new_n301), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n360), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n688), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n375), .A2(KEYINPUT101), .A3(new_n360), .A4(new_n376), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n317), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n687), .A2(new_n534), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n675), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT34), .B(G104), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G6));
  NAND2_X1  g515(.A1(new_n524), .A2(new_n527), .ZN(new_n702));
  INV_X1    g516(.A(new_n697), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT20), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n487), .A2(new_n704), .A3(new_n488), .A4(new_n489), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n495), .B1(new_n676), .B2(new_n705), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n702), .A2(new_n703), .A3(new_n535), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n675), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT35), .B(G107), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G9));
  NOR2_X1   g524(.A1(new_n628), .A2(KEYINPUT36), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n627), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n301), .A3(new_n646), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n656), .B2(new_n657), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n659), .B1(new_n593), .B2(new_n301), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n594), .B2(new_n593), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n385), .A2(new_n714), .A3(new_n537), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT37), .B(G110), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G12));
  AOI21_X1  g533(.A(new_n314), .B1(new_n645), .B2(new_n713), .ZN(new_n720));
  INV_X1    g534(.A(G900), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n529), .B1(new_n533), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n706), .A2(new_n702), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n724), .A3(new_n601), .A4(new_n703), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G128), .ZN(G30));
  INV_X1    g540(.A(new_n314), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n722), .B(KEYINPUT39), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT40), .Z(new_n730));
  XOR2_X1   g544(.A(new_n383), .B(KEYINPUT38), .Z(new_n731));
  NOR2_X1   g545(.A1(new_n491), .A2(new_n495), .ZN(new_n732));
  INV_X1    g546(.A(new_n702), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n316), .ZN(new_n734));
  INV_X1    g548(.A(new_n714), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n581), .A2(new_n582), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n542), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n560), .A2(new_n567), .ZN(new_n738));
  AOI21_X1  g552(.A(G902), .B1(new_n738), .B2(new_n543), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI22_X1  g554(.A1(new_n599), .A2(new_n600), .B1(new_n659), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n730), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n743), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n225), .ZN(G45));
  OAI211_X1 g560(.A(new_n686), .B(new_n723), .C1(new_n491), .C2(new_n495), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n720), .A2(new_n601), .A3(new_n703), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  NAND2_X1  g564(.A1(new_n299), .A2(new_n301), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n313), .A3(new_n302), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n658), .A2(new_n667), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n698), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n707), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n697), .A2(new_n753), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n714), .A2(new_n537), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n762), .B2(new_n667), .ZN(new_n763));
  INV_X1    g577(.A(new_n536), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n678), .A2(new_n679), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(G902), .B1(new_n288), .B2(new_n298), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G469), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n317), .A3(new_n313), .A4(new_n696), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT104), .A3(new_n601), .A4(new_n714), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G119), .ZN(G21));
  NOR2_X1   g586(.A1(new_n733), .A2(new_n316), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n680), .A2(new_n696), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n753), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n535), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n584), .A2(new_n592), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n566), .B2(new_n568), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n542), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n566), .A2(new_n568), .A3(new_n779), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n594), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n673), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n658), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G122), .ZN(G24));
  AOI21_X1  g602(.A(new_n785), .B1(new_n645), .B2(new_n713), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n748), .A3(new_n761), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G125), .ZN(G27));
  NAND3_X1  g605(.A1(new_n579), .A2(new_n595), .A3(new_n664), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n651), .A2(new_n645), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n310), .B(KEYINPUT106), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n302), .A2(new_n309), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n381), .A2(new_n317), .A3(new_n382), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n795), .A2(new_n796), .A3(new_n313), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n680), .A2(new_n797), .A3(new_n686), .A4(new_n723), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT42), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n671), .A2(new_n800), .A3(new_n601), .A4(new_n797), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(G131), .Z(G33));
  NAND4_X1  g617(.A1(new_n671), .A2(new_n724), .A3(new_n601), .A4(new_n797), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NAND2_X1  g619(.A1(new_n732), .A2(new_n686), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT43), .Z(new_n807));
  NOR2_X1   g621(.A1(new_n735), .A2(new_n716), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT107), .Z(new_n812));
  INV_X1    g626(.A(new_n796), .ZN(new_n813));
  INV_X1    g627(.A(new_n313), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n300), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT46), .B1(new_n818), .B2(new_n794), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n300), .B2(new_n766), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(KEYINPUT46), .A3(new_n794), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n728), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n813), .B(new_n823), .C1(new_n809), .C2(new_n810), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n812), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(new_n191), .ZN(G39));
  AND2_X1   g640(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g641(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n822), .B2(new_n828), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n748), .A2(new_n658), .A3(new_n796), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n601), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(new_n407), .ZN(G42));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n807), .A2(new_n529), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT114), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n731), .A2(new_n316), .A3(new_n775), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n786), .A3(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT50), .Z(new_n839));
  NAND2_X1  g653(.A1(new_n775), .A2(new_n796), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT116), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT117), .B1(new_n836), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n789), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n741), .A2(new_n658), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n529), .A3(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n847), .A2(new_n680), .A3(new_n686), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n836), .A2(new_n786), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n767), .A2(new_n814), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT115), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n813), .B(new_n850), .C1(new_n830), .C2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n834), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n834), .C1(new_n849), .C2(new_n853), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(G952), .B(new_n350), .C1(new_n847), .C2(new_n687), .ZN(new_n859));
  INV_X1    g673(.A(new_n850), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n761), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n843), .A2(new_n844), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT48), .ZN(new_n863));
  INV_X1    g677(.A(new_n793), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n849), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n839), .A2(KEYINPUT119), .A3(new_n845), .A4(new_n848), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n850), .A2(new_n813), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n830), .A2(new_n851), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n834), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n867), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n858), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n725), .A2(new_n749), .A3(new_n790), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n735), .A2(KEYINPUT113), .A3(new_n723), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n714), .B2(new_n722), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n774), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(new_n313), .A3(new_n741), .A4(new_n795), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n878), .B(new_n879), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n883), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT52), .B1(new_n887), .B2(new_n877), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n799), .A2(new_n801), .A3(new_n804), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n714), .A2(new_n727), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n706), .A2(new_n733), .A3(new_n723), .A4(new_n796), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(new_n667), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n785), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n748), .A2(new_n714), .A3(new_n894), .A4(new_n797), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT111), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n748), .A4(new_n797), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n763), .A2(new_n770), .B1(new_n754), .B2(new_n707), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n698), .A2(new_n754), .B1(new_n777), .B2(new_n786), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n890), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT109), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n534), .B1(new_n380), .B2(new_n384), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n651), .A2(new_n904), .A3(new_n674), .A4(new_n645), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n687), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n669), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n652), .A2(new_n668), .ZN(new_n908));
  INV_X1    g722(.A(new_n538), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n732), .A2(new_n702), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n717), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT110), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT110), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n717), .B(new_n914), .C1(new_n905), .C2(new_n911), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n910), .A2(KEYINPUT109), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n902), .A2(KEYINPUT112), .A3(new_n907), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT112), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT85), .B1(new_n671), .B2(new_n601), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n658), .A2(new_n667), .A3(new_n653), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n909), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n906), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n913), .A2(new_n915), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n907), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n890), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n889), .B1(new_n917), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n879), .B1(new_n725), .B2(new_n790), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(KEYINPUT53), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(KEYINPUT53), .B2(new_n928), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n925), .A2(new_n926), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT53), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n725), .A2(new_n790), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(KEYINPUT52), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n933), .A2(new_n886), .A3(new_n888), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n928), .B2(KEYINPUT53), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n932), .B1(KEYINPUT54), .B2(new_n938), .ZN(new_n939));
  OAI22_X1  g753(.A1(new_n876), .A2(new_n939), .B1(G952), .B2(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n731), .A2(new_n317), .A3(new_n313), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n767), .B(KEYINPUT49), .Z(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n806), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n846), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(G75));
  NOR2_X1   g759(.A1(new_n350), .A2(G952), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n938), .A2(G902), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n948), .B2(G210), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n341), .A2(new_n358), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n356), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n359), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT55), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n949), .B2(new_n953), .ZN(G51));
  XNOR2_X1  g769(.A(new_n938), .B(KEYINPUT54), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n794), .B(KEYINPUT57), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n299), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n948), .B(new_n817), .C1(new_n816), .C2(new_n815), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n946), .B1(new_n959), .B2(new_n960), .ZN(G54));
  NAND3_X1  g775(.A1(new_n948), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n487), .A2(new_n489), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n962), .A2(KEYINPUT120), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n947), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT120), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G60));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT59), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n684), .B1(new_n939), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n684), .A2(new_n969), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n946), .B(new_n970), .C1(new_n956), .C2(new_n971), .ZN(G63));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n973));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT60), .Z(new_n975));
  XOR2_X1   g789(.A(new_n712), .B(KEYINPUT121), .Z(new_n976));
  NAND3_X1  g790(.A1(new_n938), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n946), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n622), .B1(new_n640), .B2(new_n633), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n938), .B2(new_n975), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n977), .B(new_n979), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  AOI211_X1 g797(.A(KEYINPUT123), .B(new_n980), .C1(new_n938), .C2(new_n975), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n938), .A2(new_n975), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT123), .B1(new_n986), .B2(new_n980), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n977), .A2(new_n979), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n981), .A2(new_n982), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT124), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT122), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n981), .B2(new_n946), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n977), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n981), .A2(new_n992), .A3(new_n946), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n978), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n991), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(G66));
  AOI21_X1  g815(.A(new_n350), .B1(new_n531), .B2(G224), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n916), .A2(new_n907), .A3(new_n901), .A4(new_n900), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n350), .ZN(new_n1004));
  INV_X1    g818(.A(G898), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n950), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  NOR2_X1   g821(.A1(new_n580), .A2(new_n553), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n410), .A2(new_n416), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT126), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1008), .B(new_n1010), .Z(new_n1011));
  NOR2_X1   g825(.A1(new_n825), .A2(new_n832), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT62), .B1(new_n745), .B2(new_n877), .ZN(new_n1013));
  OR3_X1    g827(.A1(new_n745), .A2(KEYINPUT62), .A3(new_n877), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n687), .A2(new_n911), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n729), .A2(new_n813), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n908), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1011), .B1(new_n1018), .B2(new_n350), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n823), .A2(new_n774), .A3(new_n793), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1012), .A2(new_n878), .A3(new_n890), .A4(new_n1021), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1022), .A2(G953), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1011), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(G900), .B2(G953), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1019), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(G953), .B1(new_n188), .B2(new_n721), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1026), .B(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n1018), .B2(new_n1003), .ZN(new_n1031));
  INV_X1    g845(.A(new_n737), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1030), .B1(new_n1022), .B2(new_n1003), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n736), .A2(new_n542), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1033), .A2(new_n1036), .A3(new_n947), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1030), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n1032), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1037), .B1(new_n931), .B2(new_n1039), .ZN(G57));
endmodule


