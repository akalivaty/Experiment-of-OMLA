

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U324 ( .A1(n527), .A2(n451), .ZN(n563) );
  XOR2_X1 U325 ( .A(n422), .B(n421), .Z(n292) );
  XNOR2_X1 U326 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U327 ( .A(n397), .B(n354), .ZN(n355) );
  XNOR2_X1 U328 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U329 ( .A(n363), .B(n362), .ZN(n371) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G127GAT), .B(KEYINPUT0), .Z(n294) );
  XNOR2_X1 U334 ( .A(G113GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n318) );
  XOR2_X1 U336 ( .A(n318), .B(G120GAT), .Z(n296) );
  NAND2_X1 U337 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n311) );
  XOR2_X1 U339 ( .A(G99GAT), .B(KEYINPUT84), .Z(n298) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n301) );
  XOR2_X1 U342 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n300) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n446) );
  XOR2_X1 U345 ( .A(n301), .B(n446), .Z(n309) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n303) );
  XNOR2_X1 U347 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U349 ( .A(G176GAT), .B(G183GAT), .Z(n305) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G15GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U354 ( .A(n311), .B(n310), .Z(n527) );
  XOR2_X1 U355 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n450) );
  XOR2_X1 U356 ( .A(G120GAT), .B(G148GAT), .Z(n353) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(G85GAT), .Z(n313) );
  XNOR2_X1 U358 ( .A(G29GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U360 ( .A(n353), .B(n314), .Z(n316) );
  NAND2_X1 U361 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n317), .B(G57GAT), .Z(n320) );
  XNOR2_X1 U364 ( .A(n318), .B(KEYINPUT4), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U366 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n322) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U369 ( .A(n324), .B(n323), .Z(n333) );
  XOR2_X1 U370 ( .A(KEYINPUT2), .B(G162GAT), .Z(n326) );
  XNOR2_X1 U371 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U372 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(n327), .ZN(n349) );
  INV_X1 U374 ( .A(n349), .ZN(n331) );
  XOR2_X1 U375 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n329) );
  XNOR2_X1 U376 ( .A(KEYINPUT6), .B(KEYINPUT89), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n333), .B(n332), .ZN(n513) );
  INV_X1 U380 ( .A(n513), .ZN(n569) );
  XOR2_X1 U381 ( .A(KEYINPUT88), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(G211GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n347) );
  XOR2_X1 U384 ( .A(G155GAT), .B(G78GAT), .Z(n404) );
  XOR2_X1 U385 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n337) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U388 ( .A(n404), .B(n338), .Z(n340) );
  NAND2_X1 U389 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n341), .B(G204GAT), .Z(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n343) );
  XNOR2_X1 U393 ( .A(G197GAT), .B(G218GAT), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n436) );
  XNOR2_X1 U395 ( .A(n436), .B(KEYINPUT23), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U397 ( .A(n347), .B(n346), .Z(n348) );
  XNOR2_X1 U398 ( .A(n349), .B(n348), .ZN(n463) );
  AND2_X1 U399 ( .A1(n569), .A2(n463), .ZN(n448) );
  XOR2_X1 U400 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n351) );
  XNOR2_X1 U401 ( .A(G71GAT), .B(G57GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n397) );
  AND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT74), .B(n355), .Z(n363) );
  XOR2_X1 U405 ( .A(KEYINPUT76), .B(G85GAT), .Z(n357) );
  XNOR2_X1 U406 ( .A(G99GAT), .B(G106GAT), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n357), .B(n356), .ZN(n381) );
  XNOR2_X1 U408 ( .A(n381), .B(KEYINPUT33), .ZN(n361) );
  XOR2_X1 U409 ( .A(KEYINPUT72), .B(KEYINPUT78), .Z(n359) );
  XNOR2_X1 U410 ( .A(G78GAT), .B(KEYINPUT75), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n360) );
  XOR2_X1 U412 ( .A(G92GAT), .B(KEYINPUT79), .Z(n365) );
  XNOR2_X1 U413 ( .A(G204GAT), .B(G64GAT), .ZN(n364) );
  XNOR2_X1 U414 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U415 ( .A(G176GAT), .B(n366), .Z(n441) );
  XOR2_X1 U416 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n368) );
  XNOR2_X1 U417 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U419 ( .A(n441), .B(n369), .ZN(n370) );
  XNOR2_X1 U420 ( .A(n371), .B(n370), .ZN(n576) );
  INV_X1 U421 ( .A(n576), .ZN(n409) );
  XOR2_X1 U422 ( .A(KEYINPUT10), .B(G218GAT), .Z(n373) );
  NAND2_X1 U423 ( .A1(G232GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U425 ( .A(G92GAT), .B(G162GAT), .Z(n375) );
  XNOR2_X1 U426 ( .A(G134GAT), .B(G190GAT), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U428 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n379) );
  XNOR2_X1 U430 ( .A(KEYINPUT80), .B(KEYINPUT9), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U432 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U433 ( .A(n383), .B(n382), .ZN(n391) );
  XOR2_X1 U434 ( .A(G29GAT), .B(G36GAT), .Z(n385) );
  XNOR2_X1 U435 ( .A(G50GAT), .B(G43GAT), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U437 ( .A(KEYINPUT7), .B(KEYINPUT68), .Z(n387) );
  XNOR2_X1 U438 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U440 ( .A(n389), .B(n388), .Z(n414) );
  INV_X1 U441 ( .A(n414), .ZN(n390) );
  XOR2_X1 U442 ( .A(n391), .B(n390), .Z(n553) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(n553), .ZN(n583) );
  XOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n393) );
  NAND2_X1 U445 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U447 ( .A(n394), .B(KEYINPUT15), .Z(n399) );
  XOR2_X1 U448 ( .A(KEYINPUT69), .B(G1GAT), .Z(n396) );
  XNOR2_X1 U449 ( .A(G22GAT), .B(G15GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n415) );
  XNOR2_X1 U451 ( .A(n415), .B(n397), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT14), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U454 ( .A(G8GAT), .B(G127GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n406) );
  XOR2_X1 U457 ( .A(G183GAT), .B(G211GAT), .Z(n439) );
  XNOR2_X1 U458 ( .A(n404), .B(n439), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n482) );
  INV_X1 U460 ( .A(n482), .ZN(n579) );
  NOR2_X1 U461 ( .A1(n583), .A2(n579), .ZN(n407) );
  XOR2_X1 U462 ( .A(KEYINPUT45), .B(n407), .Z(n408) );
  NOR2_X1 U463 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U464 ( .A(KEYINPUT110), .B(n410), .ZN(n424) );
  XOR2_X1 U465 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n412) );
  XNOR2_X1 U466 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n422) );
  XOR2_X1 U469 ( .A(n415), .B(KEYINPUT30), .Z(n417) );
  NAND2_X1 U470 ( .A1(G229GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U472 ( .A(G169GAT), .B(G8GAT), .Z(n442) );
  XOR2_X1 U473 ( .A(n418), .B(n442), .Z(n420) );
  XNOR2_X1 U474 ( .A(G141GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(KEYINPUT70), .B(n292), .Z(n555) );
  INV_X1 U477 ( .A(n555), .ZN(n423) );
  NAND2_X1 U478 ( .A1(n424), .A2(n423), .ZN(n433) );
  XOR2_X1 U479 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n425) );
  XNOR2_X1 U480 ( .A(KEYINPUT47), .B(n425), .ZN(n431) );
  XOR2_X1 U481 ( .A(n482), .B(KEYINPUT106), .Z(n565) );
  XOR2_X1 U482 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n427) );
  XOR2_X1 U483 ( .A(n576), .B(KEYINPUT41), .Z(n545) );
  OR2_X1 U484 ( .A1(n292), .A2(n545), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  AND2_X1 U486 ( .A1(n565), .A2(n428), .ZN(n429) );
  AND2_X1 U487 ( .A1(n553), .A2(n429), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  AND2_X1 U489 ( .A1(n433), .A2(n432), .ZN(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n524) );
  XOR2_X1 U492 ( .A(n436), .B(G36GAT), .Z(n438) );
  NAND2_X1 U493 ( .A1(G226GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n503) );
  NOR2_X1 U499 ( .A1(n524), .A2(n503), .ZN(n447) );
  XNOR2_X1 U500 ( .A(KEYINPUT54), .B(n447), .ZN(n568) );
  NAND2_X1 U501 ( .A1(n448), .A2(n568), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U503 ( .A(n553), .ZN(n456) );
  NAND2_X1 U504 ( .A1(n563), .A2(n456), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n453) );
  XOR2_X1 U506 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n472) );
  NAND2_X1 U507 ( .A1(n576), .A2(n555), .ZN(n487) );
  NOR2_X1 U508 ( .A1(n456), .A2(n579), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT16), .ZN(n470) );
  INV_X1 U510 ( .A(n527), .ZN(n517) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n503), .Z(n461) );
  NAND2_X1 U512 ( .A1(n513), .A2(n461), .ZN(n523) );
  NOR2_X1 U513 ( .A1(n517), .A2(n523), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n463), .B(KEYINPUT28), .ZN(n525) );
  NAND2_X1 U515 ( .A1(n458), .A2(n525), .ZN(n469) );
  NOR2_X1 U516 ( .A1(n463), .A2(n517), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n570) );
  NAND2_X1 U519 ( .A1(n461), .A2(n570), .ZN(n466) );
  INV_X1 U520 ( .A(n503), .ZN(n515) );
  NAND2_X1 U521 ( .A1(n515), .A2(n517), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n569), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n484) );
  NAND2_X1 U527 ( .A1(n470), .A2(n484), .ZN(n497) );
  NOR2_X1 U528 ( .A1(n487), .A2(n497), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n479), .A2(n513), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n479), .A2(n515), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT96), .ZN(n475) );
  XNOR2_X1 U534 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U536 ( .A1(n479), .A2(n517), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U538 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  INV_X1 U539 ( .A(n525), .ZN(n519) );
  NAND2_X1 U540 ( .A1(n479), .A2(n519), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT98), .ZN(n481) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U543 ( .A1(n583), .A2(n482), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT99), .B(n486), .ZN(n511) );
  NOR2_X1 U547 ( .A1(n511), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT38), .B(n488), .ZN(n495) );
  NAND2_X1 U549 ( .A1(n513), .A2(n495), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n515), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n495), .A2(n517), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U558 ( .A1(n519), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n496), .ZN(G1331GAT) );
  INV_X1 U560 ( .A(n545), .ZN(n560) );
  NAND2_X1 U561 ( .A1(n292), .A2(n560), .ZN(n510) );
  NOR2_X1 U562 ( .A1(n510), .A2(n497), .ZN(n498) );
  XOR2_X1 U563 ( .A(KEYINPUT102), .B(n498), .Z(n506) );
  NOR2_X1 U564 ( .A1(n569), .A2(n506), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n500) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n506), .A2(n503), .ZN(n504) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n527), .A2(n506), .ZN(n505) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n506), .A2(n525), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U578 ( .A(KEYINPUT105), .B(n512), .Z(n520) );
  NAND2_X1 U579 ( .A1(n513), .A2(n520), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n520), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n520), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n540) );
  NAND2_X1 U589 ( .A1(n540), .A2(n525), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n555), .A2(n531), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n560), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  INV_X1 U596 ( .A(n531), .ZN(n535) );
  NOR2_X1 U597 ( .A1(n565), .A2(n535), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U601 ( .A1(n535), .A2(n553), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n537) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n570), .A2(n540), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n292), .A2(n552), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n549) );
  NOR2_X1 U613 ( .A1(n545), .A2(n552), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n579), .A2(n552), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n563), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(n559), .Z(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  INV_X1 U630 ( .A(n563), .ZN(n564) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  AND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n582) );
  NOR2_X1 U636 ( .A1(n582), .A2(n292), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n582), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n582), .ZN(n580) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(n580), .Z(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

