//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(G43gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT15), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n207), .B1(new_n213), .B2(KEYINPUT82), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT82), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n203), .B(KEYINPUT84), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n204), .B(KEYINPUT83), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT15), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n207), .B(KEYINPUT85), .Z(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(new_n205), .A3(new_n213), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n216), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G8gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n222), .B(KEYINPUT17), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n222), .B(new_n227), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n232), .B(KEYINPUT13), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G197gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT11), .B(G169gat), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT12), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT18), .B1(new_n231), .B2(new_n232), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n243), .B1(new_n237), .B2(new_n245), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G169gat), .ZN(new_n255));
  INV_X1    g054(.A(G176gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT23), .ZN(new_n260));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT25), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT24), .ZN(new_n264));
  INV_X1    g063(.A(G183gat), .ZN(new_n265));
  INV_X1    g064(.A(G190gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n268));
  MUX2_X1   g067(.A(G183gat), .B(new_n268), .S(G190gat), .Z(new_n269));
  AOI21_X1  g068(.A(new_n263), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n271), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT25), .B1(new_n274), .B2(new_n262), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n266), .ZN(new_n279));
  INV_X1    g078(.A(new_n277), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT28), .B1(new_n280), .B2(G190gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n257), .A2(new_n282), .A3(new_n261), .ZN(new_n283));
  OAI221_X1 g082(.A(new_n283), .B1(new_n282), .B2(new_n257), .C1(new_n265), .C2(new_n266), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n279), .B(new_n281), .C1(new_n284), .C2(KEYINPUT65), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n254), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n253), .B1(new_n276), .B2(new_n287), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G211gat), .B(G218gat), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT67), .B(G197gat), .ZN(new_n295));
  INV_X1    g094(.A(G204gat), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI22_X1  g100(.A1(new_n297), .A2(new_n298), .B1(KEYINPUT22), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(new_n293), .A3(new_n303), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n288), .A2(new_n254), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n276), .B2(new_n287), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(new_n254), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n317), .B1(new_n320), .B2(KEYINPUT69), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n310), .B(new_n316), .C1(new_n321), .C2(new_n309), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT72), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT69), .B1(new_n290), .B2(new_n291), .ZN(new_n325));
  INV_X1    g124(.A(new_n317), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n309), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n310), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n315), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n323), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n324), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n334));
  XOR2_X1   g133(.A(G1gat), .B(G29gat), .Z(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G57gat), .B(G85gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G127gat), .B(G134gat), .Z(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  XOR2_X1   g140(.A(G113gat), .B(G120gat), .Z(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n343), .B(new_n345), .Z(new_n346));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  OR2_X1    g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(KEYINPUT2), .ZN(new_n349));
  INV_X1    g148(.A(G141gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G148gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(G148gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(KEYINPUT73), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n354), .A2(new_n350), .A3(G148gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G141gat), .B(G148gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n347), .B(new_n348), .C1(new_n357), .C2(KEYINPUT2), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n359), .B(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(new_n346), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n343), .B(new_n345), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n360), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n366), .B(new_n370), .C1(KEYINPUT4), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n359), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n365), .B1(new_n375), .B2(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n365), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n371), .A2(new_n360), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n373), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT75), .B1(new_n382), .B2(KEYINPUT5), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n374), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n359), .B(KEYINPUT74), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n371), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n387), .B(KEYINPUT77), .C1(new_n386), .C2(new_n373), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n378), .A4(new_n366), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n334), .B(new_n339), .C1(new_n384), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n339), .A3(new_n390), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n339), .B1(new_n384), .B2(new_n390), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n334), .B(new_n393), .C1(new_n394), .C2(KEYINPUT78), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n320), .A2(new_n328), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n327), .B2(new_n328), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT72), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT30), .A4(new_n316), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n333), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n306), .A2(new_n308), .A3(new_n289), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT3), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT79), .A4(new_n289), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n360), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n309), .B1(new_n289), .B2(new_n362), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n385), .B1(new_n407), .B2(new_n361), .ZN(new_n414));
  OR3_X1    g213(.A1(new_n412), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n413), .B2(new_n415), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n405), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G15gat), .B(G43gat), .Z(new_n422));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n276), .A2(new_n346), .A3(new_n287), .ZN(new_n426));
  INV_X1    g225(.A(G227gat), .ZN(new_n427));
  INV_X1    g226(.A(G233gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n270), .A2(new_n275), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n285), .A2(new_n286), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n371), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n425), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n426), .A2(new_n432), .ZN(new_n437));
  INV_X1    g236(.A(new_n429), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT34), .B(new_n429), .C1(new_n426), .C2(new_n432), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n433), .A2(KEYINPUT32), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n437), .A2(new_n438), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT34), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n447), .B(new_n449), .C1(new_n450), .C2(new_n425), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n446), .B1(new_n451), .B2(new_n441), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n413), .A2(new_n415), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n416), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n404), .A3(new_n418), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n421), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n402), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n324), .A2(new_n331), .A3(new_n401), .A4(new_n332), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n393), .A2(new_n334), .ZN(new_n462));
  INV_X1    g261(.A(new_n394), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n391), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n421), .A2(new_n456), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n421), .A2(KEYINPUT80), .A3(new_n456), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n402), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n468), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n310), .C1(new_n321), .C2(new_n309), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n315), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n329), .B2(new_n310), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n292), .B2(new_n328), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n321), .B2(new_n328), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n475), .A2(new_n480), .A3(new_n481), .A4(new_n315), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n464), .A2(new_n478), .A3(new_n322), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n375), .A2(new_n365), .A3(new_n372), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT81), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n388), .A2(new_n389), .A3(new_n364), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n380), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n491), .A3(new_n380), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n490), .A2(KEYINPUT40), .A3(new_n339), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n463), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n492), .A2(new_n339), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT40), .B1(new_n495), .B2(new_n490), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n460), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n473), .A2(new_n483), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n445), .B2(new_n452), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n444), .B1(new_n442), .B2(new_n443), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n451), .A2(new_n446), .A3(new_n441), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n472), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n252), .B1(new_n467), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  INV_X1    g307(.A(G85gat), .ZN(new_n509));
  INV_X1    g308(.A(G92gat), .ZN(new_n510));
  AOI22_X1  g309(.A1(KEYINPUT8), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT7), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT92), .ZN(new_n515));
  AND2_X1   g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT92), .B(new_n514), .C1(new_n509), .C2(new_n510), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT93), .B1(new_n517), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G99gat), .B(G106gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n522), .B(new_n511), .C1(new_n519), .C2(new_n520), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT94), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(KEYINPUT94), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n229), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(new_n518), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n522), .B1(new_n534), .B2(new_n511), .ZN(new_n535));
  INV_X1    g334(.A(new_n525), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n537), .A2(new_n222), .B1(KEYINPUT41), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n529), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G190gat), .B(G218gat), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n538), .A2(KEYINPUT41), .ZN(new_n544));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n543), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n557), .A2(new_n555), .ZN(new_n560));
  INV_X1    g359(.A(G64gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G57gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT88), .B(G57gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n535), .B2(new_n536), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n556), .A2(new_n558), .B1(new_n564), .B2(new_n560), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n524), .A2(new_n569), .A3(new_n525), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n537), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n570), .ZN(new_n579));
  INV_X1    g378(.A(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT95), .Z(new_n583));
  AOI21_X1  g382(.A(KEYINPUT96), .B1(new_n573), .B2(new_n574), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n585));
  AOI211_X1 g384(.A(new_n585), .B(new_n580), .C1(new_n571), .C2(new_n572), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n581), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n227), .B1(KEYINPUT21), .B2(new_n569), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT89), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT91), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n548), .A2(new_n590), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n507), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n397), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(G1gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(G1324gat));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  INV_X1    g412(.A(new_n460), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT16), .B(G8gat), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G8gat), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n608), .B2(new_n460), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT42), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(KEYINPUT42), .B2(new_n616), .ZN(G1325gat));
  AND3_X1   g419(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT98), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT98), .B1(new_n501), .B2(new_n504), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(G15gat), .B1(new_n613), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n453), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n625), .A2(G15gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n613), .B2(new_n626), .ZN(G1326gat));
  NAND2_X1  g426(.A1(new_n470), .A2(new_n471), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n608), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT43), .B(G22gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1327gat));
  INV_X1    g431(.A(new_n606), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n590), .A2(new_n547), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n507), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n208), .A3(new_n609), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT45), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n458), .A2(KEYINPUT35), .B1(new_n461), .B2(new_n465), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n472), .A2(new_n499), .A3(new_n623), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n472), .A2(new_n623), .A3(new_n499), .A4(KEYINPUT101), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n639), .B1(new_n645), .B2(new_n547), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n467), .A2(new_n506), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(KEYINPUT44), .A3(new_n548), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n606), .B(KEYINPUT99), .ZN(new_n650));
  INV_X1    g449(.A(new_n590), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n251), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT100), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G29gat), .B1(new_n654), .B2(new_n397), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n655), .ZN(G1328gat));
  NOR3_X1   g455(.A1(new_n635), .A2(G36gat), .A3(new_n614), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT46), .ZN(new_n658));
  INV_X1    g457(.A(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n460), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT102), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(G36gat), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(KEYINPUT102), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(G1329gat));
  AOI21_X1  g463(.A(G43gat), .B1(new_n636), .B2(new_n453), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(KEYINPUT103), .B2(KEYINPUT47), .ZN(new_n666));
  INV_X1    g465(.A(new_n623), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G43gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n654), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(G1330gat));
  OAI21_X1  g470(.A(G50gat), .B1(new_n654), .B2(new_n473), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n635), .A2(G50gat), .A3(new_n628), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(KEYINPUT48), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n629), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n676), .B2(G50gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g477(.A1(new_n547), .A2(new_n633), .ZN(new_n679));
  NOR4_X1   g478(.A1(new_n645), .A2(new_n251), .A3(new_n679), .A4(new_n651), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n397), .B(KEYINPUT104), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT105), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n563), .ZN(G1332gat));
  AOI21_X1  g484(.A(new_n614), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT106), .Z(new_n688));
  NOR2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1333gat));
  AOI21_X1  g489(.A(new_n553), .B1(new_n680), .B2(new_n667), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n625), .A2(G71gat), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n680), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g493(.A1(new_n680), .A2(new_n629), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(G78gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1335gat));
  NOR2_X1   g496(.A1(new_n633), .A2(new_n251), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n651), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n649), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G85gat), .B1(new_n702), .B2(new_n397), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n643), .A2(new_n644), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n548), .B(new_n698), .C1(new_n704), .C2(new_n640), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n645), .A2(new_n547), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n698), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n651), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n509), .A3(new_n609), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(new_n711), .ZN(G1336gat));
  NAND2_X1  g511(.A1(new_n701), .A2(new_n460), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n707), .A2(new_n709), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n460), .A2(new_n510), .A3(new_n590), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT108), .Z(new_n716));
  AOI22_X1  g515(.A1(new_n713), .A2(G92gat), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1337gat));
  OAI21_X1  g518(.A(G99gat), .B1(new_n702), .B2(new_n623), .ZN(new_n720));
  INV_X1    g519(.A(G99gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n710), .A2(new_n721), .A3(new_n453), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1338gat));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n473), .A2(G106gat), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n646), .A2(new_n629), .A3(new_n648), .A4(new_n700), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G106gat), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n710), .A2(new_n725), .B1(new_n727), .B2(KEYINPUT109), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n729), .A3(G106gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n724), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n649), .A2(new_n468), .A3(new_n700), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G106gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n710), .A2(new_n725), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT111), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n738), .A3(new_n730), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT53), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n737), .A2(new_n743), .ZN(G1339gat));
  NAND2_X1  g543(.A1(new_n607), .A2(new_n252), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n582), .B(KEYINPUT95), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n573), .A2(new_n574), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n580), .B1(new_n571), .B2(new_n572), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n584), .A2(new_n586), .A3(KEYINPUT54), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT112), .B1(new_n751), .B2(new_n578), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n575), .A2(new_n585), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(KEYINPUT96), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n748), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n588), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n750), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n746), .B1(new_n758), .B2(KEYINPUT55), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n234), .A2(new_n235), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT113), .Z(new_n761));
  NOR2_X1   g560(.A1(new_n231), .A2(new_n232), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n241), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n249), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n547), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n750), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n751), .A2(KEYINPUT112), .A3(new_n578), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n756), .B1(new_n755), .B2(new_n588), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n759), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n764), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n590), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n251), .B1(new_n758), .B2(KEYINPUT55), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT55), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n583), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n772), .B1(new_n547), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n650), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n745), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n682), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(new_n460), .A3(new_n457), .ZN(new_n783));
  AOI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n251), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n628), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n614), .A2(new_n609), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n785), .A2(new_n625), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n251), .A2(G113gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(G1340gat));
  AOI21_X1  g588(.A(G120gat), .B1(new_n783), .B2(new_n590), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n590), .A2(G120gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n787), .B2(new_n791), .ZN(G1341gat));
  INV_X1    g591(.A(new_n787), .ZN(new_n793));
  OAI21_X1  g592(.A(G127gat), .B1(new_n793), .B2(new_n650), .ZN(new_n794));
  INV_X1    g593(.A(G127gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n795), .A3(new_n633), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1342gat));
  INV_X1    g596(.A(G134gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n798), .A3(new_n548), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n799), .A2(KEYINPUT56), .ZN(new_n800));
  OAI21_X1  g599(.A(G134gat), .B1(new_n793), .B2(new_n547), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(KEYINPUT56), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(G1343gat));
  NOR2_X1   g602(.A1(new_n667), .A2(new_n786), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n548), .B1(new_n778), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n774), .B(KEYINPUT116), .C1(new_n775), .C2(new_n777), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n772), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n810), .B2(new_n809), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n606), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n745), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT57), .A3(new_n629), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n781), .A2(new_n468), .ZN(new_n816));
  XOR2_X1   g615(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n805), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n251), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G141gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824));
  INV_X1    g623(.A(new_n782), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n667), .A2(new_n460), .A3(new_n473), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(G141gat), .A3(new_n252), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n823), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n350), .B1(new_n821), .B2(new_n251), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT58), .B1(new_n831), .B2(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  INV_X1    g632(.A(new_n827), .ZN(new_n834));
  INV_X1    g633(.A(G148gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n590), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n745), .B(KEYINPUT118), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n772), .B1(new_n807), .B2(new_n808), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n633), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n628), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n837), .B(KEYINPUT119), .C1(new_n838), .C2(new_n633), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT57), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n816), .A2(new_n817), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n845), .A2(new_n651), .A3(new_n667), .A4(new_n786), .ZN(new_n846));
  NAND2_X1  g645(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n835), .B1(new_n821), .B2(new_n590), .ZN(new_n848));
  OAI221_X1 g647(.A(new_n836), .B1(new_n846), .B2(new_n847), .C1(new_n848), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g648(.A(G155gat), .B1(new_n834), .B2(new_n633), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n780), .A2(G155gat), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT120), .Z(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n821), .B2(new_n852), .ZN(G1346gat));
  AOI21_X1  g652(.A(G162gat), .B1(new_n834), .B2(new_n548), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n548), .A2(G162gat), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n821), .B2(new_n855), .ZN(G1347gat));
  NAND2_X1  g655(.A1(new_n681), .A2(new_n460), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n625), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT122), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n628), .A3(new_n781), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n255), .A3(new_n252), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n781), .A2(new_n397), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n460), .A3(new_n473), .A4(new_n453), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT121), .Z(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n251), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n865), .B2(new_n255), .ZN(G1348gat));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n256), .A3(new_n590), .ZN(new_n867));
  OAI21_X1  g666(.A(G176gat), .B1(new_n860), .B2(new_n651), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1349gat));
  OAI21_X1  g668(.A(G183gat), .B1(new_n860), .B2(new_n650), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n633), .A2(new_n277), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(KEYINPUT123), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n872), .B(new_n874), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n864), .A2(new_n266), .A3(new_n548), .ZN(new_n876));
  OAI21_X1  g675(.A(G190gat), .B1(new_n860), .B2(new_n547), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT61), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1351gat));
  AND4_X1   g678(.A1(new_n460), .A2(new_n862), .A3(new_n468), .A4(new_n623), .ZN(new_n880));
  XOR2_X1   g679(.A(KEYINPUT124), .B(G197gat), .Z(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n251), .A3(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT125), .Z(new_n883));
  NOR2_X1   g682(.A1(new_n857), .A2(new_n667), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n843), .B2(new_n844), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n252), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n886), .B2(new_n881), .ZN(G1352gat));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n296), .A3(new_n590), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT62), .Z(new_n889));
  NOR2_X1   g688(.A1(new_n885), .A2(new_n651), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n889), .B(KEYINPUT126), .C1(new_n296), .C2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(new_n296), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n888), .B(KEYINPUT62), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n891), .A2(new_n895), .ZN(G1353gat));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n299), .A3(new_n633), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n633), .B(new_n884), .C1(new_n843), .C2(new_n844), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n898), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT63), .B1(new_n898), .B2(G211gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT127), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1354gat));
  OAI21_X1  g704(.A(G218gat), .B1(new_n885), .B2(new_n547), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n880), .A2(new_n300), .A3(new_n548), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1355gat));
endmodule


