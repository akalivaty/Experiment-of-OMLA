

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G2105), .A2(n517), .ZN(n886) );
  NOR2_X1 U555 ( .A1(n691), .A2(n690), .ZN(n693) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n692) );
  NOR2_X1 U557 ( .A1(n526), .A2(n525), .ZN(G160) );
  OR2_X1 U558 ( .A1(n777), .A2(n766), .ZN(n516) );
  NOR2_X1 U559 ( .A1(n746), .A2(n748), .ZN(n682) );
  INV_X1 U560 ( .A(KEYINPUT102), .ZN(n715) );
  NOR2_X1 U561 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U562 ( .A(KEYINPUT103), .B(KEYINPUT29), .ZN(n724) );
  XNOR2_X1 U563 ( .A(n725), .B(n724), .ZN(n728) );
  NOR2_X1 U564 ( .A1(G1384), .A2(G164), .ZN(n678) );
  NAND2_X1 U565 ( .A1(n516), .A2(n1010), .ZN(n767) );
  NOR2_X1 U566 ( .A1(G651), .A2(n629), .ZN(n649) );
  AND2_X1 U567 ( .A1(n533), .A2(n532), .ZN(G164) );
  INV_X1 U568 ( .A(G2104), .ZN(n517) );
  INV_X1 U569 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U570 ( .A1(n517), .A2(n522), .ZN(n527) );
  NAND2_X1 U571 ( .A1(n527), .A2(G113), .ZN(n520) );
  NAND2_X1 U572 ( .A1(G101), .A2(n886), .ZN(n518) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U574 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n521), .Z(n887) );
  NAND2_X1 U577 ( .A1(G137), .A2(n887), .ZN(n524) );
  NOR2_X1 U578 ( .A1(n522), .A2(G2104), .ZN(n890) );
  NAND2_X1 U579 ( .A1(G125), .A2(n890), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n887), .A2(G138), .ZN(n533) );
  AND2_X1 U582 ( .A1(G114), .A2(n527), .ZN(n529) );
  AND2_X1 U583 ( .A1(G126), .A2(n890), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G102), .A2(n886), .ZN(n530) );
  AND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U587 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U588 ( .A1(G123), .A2(n890), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n534), .B(KEYINPUT18), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G99), .A2(n886), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G135), .A2(n887), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n527), .A2(G111), .ZN(n537) );
  XOR2_X1 U594 ( .A(KEYINPUT82), .B(n537), .Z(n538) );
  NOR2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n940) );
  XNOR2_X1 U597 ( .A(G2096), .B(n940), .ZN(n542) );
  OR2_X1 U598 ( .A1(G2100), .A2(n542), .ZN(G156) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  XNOR2_X1 U600 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n549) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n543) );
  XOR2_X1 U602 ( .A(KEYINPUT65), .B(n543), .Z(n643) );
  NAND2_X1 U603 ( .A1(G90), .A2(n643), .ZN(n546) );
  INV_X1 U604 ( .A(G651), .ZN(n551) );
  XOR2_X1 U605 ( .A(G543), .B(KEYINPUT0), .Z(n544) );
  XNOR2_X1 U606 ( .A(KEYINPUT66), .B(n544), .ZN(n629) );
  NOR2_X1 U607 ( .A1(n551), .A2(n629), .ZN(n639) );
  NAND2_X1 U608 ( .A1(G77), .A2(n639), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT9), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n549), .B(n548), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n649), .A2(G52), .ZN(n550) );
  XNOR2_X1 U613 ( .A(n550), .B(KEYINPUT68), .ZN(n554) );
  NOR2_X1 U614 ( .A1(G543), .A2(n551), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT1), .B(n552), .Z(n642) );
  NAND2_X1 U616 ( .A1(G64), .A2(n642), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(G88), .A2(n643), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G75), .A2(n639), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G62), .A2(n642), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G50), .A2(n649), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G65), .A2(n642), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G78), .A2(n639), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G91), .A2(n643), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT71), .B(n565), .ZN(n566) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n649), .A2(G53), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(G299) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT74), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT10), .B(n571), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n832) );
  NAND2_X1 U639 ( .A1(n832), .A2(G567), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  NAND2_X1 U641 ( .A1(n643), .A2(G81), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G68), .A2(n639), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n576), .Z(n580) );
  NAND2_X1 U646 ( .A1(G56), .A2(n642), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT14), .ZN(n578) );
  XNOR2_X1 U648 ( .A(n578), .B(KEYINPUT75), .ZN(n579) );
  NOR2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n649), .A2(G43), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n995) );
  INV_X1 U652 ( .A(G860), .ZN(n609) );
  OR2_X1 U653 ( .A1(n995), .A2(n609), .ZN(G153) );
  NAND2_X1 U654 ( .A1(G301), .A2(G868), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT76), .ZN(n594) );
  INV_X1 U656 ( .A(G868), .ZN(n661) );
  NAND2_X1 U657 ( .A1(n643), .A2(G92), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G54), .A2(n649), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G79), .A2(n639), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U661 ( .A(KEYINPUT78), .B(n586), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G66), .A2(n642), .ZN(n587) );
  XNOR2_X1 U663 ( .A(KEYINPUT77), .B(n587), .ZN(n588) );
  NOR2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n592), .Z(n610) );
  NAND2_X1 U667 ( .A1(n661), .A2(n610), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U669 ( .A1(n643), .A2(G89), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n595), .B(KEYINPUT4), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G76), .A2(n639), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT5), .ZN(n604) );
  XNOR2_X1 U674 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G63), .A2(n642), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G51), .A2(n649), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U678 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT7), .B(n605), .ZN(G168) );
  XOR2_X1 U681 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(KEYINPUT80), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n661), .A2(G286), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n609), .A2(G559), .ZN(n611) );
  INV_X1 U687 ( .A(n610), .ZN(n992) );
  NAND2_X1 U688 ( .A1(n611), .A2(n992), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n995), .ZN(n613) );
  XOR2_X1 U691 ( .A(KEYINPUT81), .B(n613), .Z(n616) );
  NAND2_X1 U692 ( .A1(G868), .A2(n992), .ZN(n614) );
  NOR2_X1 U693 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G93), .A2(n643), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G80), .A2(n639), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G67), .A2(n642), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G55), .A2(n649), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n660) );
  NAND2_X1 U702 ( .A1(n992), .A2(G559), .ZN(n658) );
  XOR2_X1 U703 ( .A(KEYINPUT83), .B(n995), .Z(n623) );
  XNOR2_X1 U704 ( .A(n658), .B(n623), .ZN(n624) );
  NOR2_X1 U705 ( .A1(G860), .A2(n624), .ZN(n625) );
  XOR2_X1 U706 ( .A(n660), .B(n625), .Z(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n649), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n642), .A2(n628), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G87), .A2(n629), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U713 ( .A1(n649), .A2(G47), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n642), .A2(G60), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U716 ( .A(KEYINPUT67), .B(n634), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G85), .A2(n643), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G72), .A2(n639), .ZN(n635) );
  AND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G290) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n641) );
  NAND2_X1 U722 ( .A1(G73), .A2(n639), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n641), .B(n640), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G61), .A2(n642), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G86), .A2(n643), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U728 ( .A(KEYINPUT85), .B(n648), .Z(n651) );
  NAND2_X1 U729 ( .A1(n649), .A2(G48), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G305) );
  XNOR2_X1 U731 ( .A(n660), .B(KEYINPUT19), .ZN(n652) );
  XNOR2_X1 U732 ( .A(G288), .B(n652), .ZN(n655) );
  XNOR2_X1 U733 ( .A(G166), .B(G290), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(G299), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(G305), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n995), .B(n657), .ZN(n900) );
  XNOR2_X1 U738 ( .A(n658), .B(n900), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT86), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(G2072), .A2(n668), .ZN(G158) );
  XOR2_X1 U748 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U749 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U751 ( .A1(G120), .A2(G108), .ZN(n669) );
  NOR2_X1 U752 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(G69), .A2(n670), .ZN(n836) );
  NAND2_X1 U754 ( .A1(n836), .A2(G567), .ZN(n676) );
  NOR2_X1 U755 ( .A1(G219), .A2(G220), .ZN(n672) );
  XNOR2_X1 U756 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n671) );
  XNOR2_X1 U757 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U758 ( .A1(n673), .A2(G218), .ZN(n674) );
  NAND2_X1 U759 ( .A1(G96), .A2(n674), .ZN(n837) );
  NAND2_X1 U760 ( .A1(n837), .A2(G2106), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n838) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U763 ( .A1(n838), .A2(n677), .ZN(n835) );
  NAND2_X1 U764 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n782) );
  INV_X1 U767 ( .A(n782), .ZN(n679) );
  XNOR2_X1 U768 ( .A(n678), .B(KEYINPUT64), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n679), .A2(n708), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G8), .A2(n681), .ZN(n731) );
  NOR2_X1 U771 ( .A1(G1966), .A2(n731), .ZN(n680) );
  XOR2_X1 U772 ( .A(KEYINPUT95), .B(n680), .Z(n746) );
  INV_X1 U773 ( .A(n681), .ZN(n707) );
  INV_X1 U774 ( .A(n707), .ZN(n733) );
  NOR2_X1 U775 ( .A1(G2084), .A2(n733), .ZN(n748) );
  NAND2_X1 U776 ( .A1(G8), .A2(n682), .ZN(n683) );
  XNOR2_X1 U777 ( .A(KEYINPUT30), .B(n683), .ZN(n684) );
  XNOR2_X1 U778 ( .A(n684), .B(KEYINPUT104), .ZN(n685) );
  NOR2_X1 U779 ( .A1(n685), .A2(G168), .ZN(n691) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .ZN(n927) );
  NAND2_X1 U781 ( .A1(n707), .A2(n927), .ZN(n686) );
  XOR2_X1 U782 ( .A(KEYINPUT96), .B(n686), .Z(n688) );
  NOR2_X1 U783 ( .A1(n707), .A2(G1961), .ZN(n687) );
  XNOR2_X1 U784 ( .A(KEYINPUT97), .B(n689), .ZN(n726) );
  NOR2_X1 U785 ( .A1(G171), .A2(n726), .ZN(n690) );
  XNOR2_X1 U786 ( .A(n693), .B(n692), .ZN(n730) );
  INV_X1 U787 ( .A(G1348), .ZN(n979) );
  NOR2_X1 U788 ( .A1(n707), .A2(n979), .ZN(n694) );
  XNOR2_X1 U789 ( .A(n694), .B(KEYINPUT101), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n707), .A2(G2067), .ZN(n695) );
  NAND2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n702) );
  INV_X1 U792 ( .A(G1996), .ZN(n920) );
  NOR2_X1 U793 ( .A1(n733), .A2(n920), .ZN(n697) );
  XOR2_X1 U794 ( .A(KEYINPUT26), .B(n697), .Z(n700) );
  AND2_X1 U795 ( .A1(n733), .A2(G1341), .ZN(n698) );
  NOR2_X1 U796 ( .A1(n698), .A2(n995), .ZN(n699) );
  AND2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n703), .A2(n992), .ZN(n701) );
  NAND2_X1 U799 ( .A1(n702), .A2(n701), .ZN(n705) );
  OR2_X1 U800 ( .A1(n703), .A2(n992), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n718) );
  INV_X1 U802 ( .A(G1956), .ZN(n706) );
  OR2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n713) );
  INV_X1 U804 ( .A(G2072), .ZN(n953) );
  NOR2_X1 U805 ( .A1(n782), .A2(n953), .ZN(n709) );
  AND2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U807 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n710) );
  XNOR2_X1 U808 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U810 ( .A(KEYINPUT99), .B(n714), .Z(n719) );
  NOR2_X1 U811 ( .A1(G299), .A2(n719), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n718), .A2(n717), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n719), .A2(G299), .ZN(n720) );
  XNOR2_X1 U815 ( .A(n720), .B(KEYINPUT28), .ZN(n721) );
  XNOR2_X1 U816 ( .A(n721), .B(KEYINPUT100), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G171), .A2(n726), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n744) );
  NAND2_X1 U821 ( .A1(n744), .A2(G286), .ZN(n739) );
  INV_X1 U822 ( .A(n731), .ZN(n732) );
  INV_X1 U823 ( .A(n732), .ZN(n777) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n777), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n736), .A2(G303), .ZN(n737) );
  XOR2_X1 U828 ( .A(KEYINPUT107), .B(n737), .Z(n738) );
  NAND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U831 ( .A(n741), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  AND2_X1 U833 ( .A1(n770), .A2(n1004), .ZN(n743) );
  INV_X1 U834 ( .A(KEYINPUT108), .ZN(n762) );
  OR2_X1 U835 ( .A1(n777), .A2(n762), .ZN(n757) );
  INV_X1 U836 ( .A(n757), .ZN(n742) );
  AND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n752) );
  XNOR2_X1 U838 ( .A(KEYINPUT105), .B(n744), .ZN(n745) );
  NOR2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U840 ( .A(KEYINPUT106), .B(n747), .ZN(n751) );
  NAND2_X1 U841 ( .A1(G8), .A2(n748), .ZN(n749) );
  XNOR2_X1 U842 ( .A(KEYINPUT94), .B(n749), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n769) );
  AND2_X1 U844 ( .A1(n752), .A2(n769), .ZN(n761) );
  INV_X1 U845 ( .A(n1004), .ZN(n755) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  NOR2_X1 U848 ( .A1(n753), .A2(n1002), .ZN(n754) );
  OR2_X1 U849 ( .A1(n755), .A2(n754), .ZN(n756) );
  OR2_X1 U850 ( .A1(n757), .A2(n756), .ZN(n759) );
  INV_X1 U851 ( .A(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U853 ( .A1(n761), .A2(n760), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n762), .A2(n1002), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n1002), .A2(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n763), .A2(KEYINPUT108), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n1010) );
  NOR2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n781) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U862 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n774), .A2(n777), .ZN(n779) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U866 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  OR2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n806) );
  XNOR2_X1 U870 ( .A(G1986), .B(G290), .ZN(n997) );
  NOR2_X1 U871 ( .A1(n782), .A2(n708), .ZN(n826) );
  NAND2_X1 U872 ( .A1(n997), .A2(n826), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(KEYINPUT88), .ZN(n804) );
  NAND2_X1 U874 ( .A1(G107), .A2(n527), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G131), .A2(n887), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G95), .A2(n886), .ZN(n786) );
  XNOR2_X1 U878 ( .A(KEYINPUT89), .B(n786), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n890), .A2(G119), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n867) );
  XNOR2_X1 U882 ( .A(KEYINPUT90), .B(G1991), .ZN(n923) );
  NAND2_X1 U883 ( .A1(n867), .A2(n923), .ZN(n802) );
  NAND2_X1 U884 ( .A1(n527), .A2(G117), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT91), .B(n791), .Z(n793) );
  NAND2_X1 U886 ( .A1(n890), .A2(G129), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U888 ( .A(KEYINPUT92), .B(n794), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G105), .A2(n886), .ZN(n795) );
  XNOR2_X1 U890 ( .A(n795), .B(KEYINPUT93), .ZN(n796) );
  XNOR2_X1 U891 ( .A(n796), .B(KEYINPUT38), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n887), .A2(G141), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n869) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n869), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n946) );
  NAND2_X1 U897 ( .A1(n946), .A2(n826), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n816) );
  XNOR2_X1 U900 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NAND2_X1 U901 ( .A1(G104), .A2(n886), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G140), .A2(n887), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U904 ( .A(KEYINPUT34), .B(n809), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G116), .A2(n527), .ZN(n811) );
  NAND2_X1 U906 ( .A1(G128), .A2(n890), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U908 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U910 ( .A(KEYINPUT36), .B(n815), .ZN(n896) );
  NOR2_X1 U911 ( .A1(n824), .A2(n896), .ZN(n949) );
  NAND2_X1 U912 ( .A1(n826), .A2(n949), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n816), .A2(n823), .ZN(n830) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n869), .ZN(n958) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n923), .A2(n867), .ZN(n942) );
  NOR2_X1 U917 ( .A1(n817), .A2(n942), .ZN(n818) );
  NOR2_X1 U918 ( .A1(n946), .A2(n818), .ZN(n819) );
  NOR2_X1 U919 ( .A1(n958), .A2(n819), .ZN(n820) );
  XOR2_X1 U920 ( .A(n820), .B(KEYINPUT39), .Z(n821) );
  XNOR2_X1 U921 ( .A(KEYINPUT109), .B(n821), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n824), .A2(n896), .ZN(n947) );
  NAND2_X1 U924 ( .A1(n825), .A2(n947), .ZN(n827) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n828), .B(KEYINPUT110), .ZN(n829) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U931 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G188) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(G325) );
  XOR2_X1 U935 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  XNOR2_X1 U936 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  INV_X1 U941 ( .A(n838), .ZN(G319) );
  XOR2_X1 U942 ( .A(KEYINPUT113), .B(G2090), .Z(n840) );
  XNOR2_X1 U943 ( .A(G2072), .B(G2078), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U945 ( .A(n841), .B(G2100), .Z(n843) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2084), .ZN(n842) );
  XNOR2_X1 U947 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U948 ( .A(G2096), .B(G2678), .Z(n845) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U950 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U951 ( .A(n847), .B(n846), .Z(G227) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1976), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1991), .B(G1996), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n850), .B(KEYINPUT114), .Z(n852) );
  XNOR2_X1 U956 ( .A(G1966), .B(G1956), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U958 ( .A(G1981), .B(G1971), .Z(n854) );
  XNOR2_X1 U959 ( .A(G1986), .B(G1961), .ZN(n853) );
  XNOR2_X1 U960 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U961 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U962 ( .A(KEYINPUT115), .B(G2474), .ZN(n857) );
  XNOR2_X1 U963 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G100), .A2(n886), .ZN(n860) );
  NAND2_X1 U965 ( .A1(G112), .A2(n527), .ZN(n859) );
  NAND2_X1 U966 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U968 ( .A(n861), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G136), .A2(n887), .ZN(n862) );
  XNOR2_X1 U970 ( .A(n862), .B(KEYINPUT116), .ZN(n863) );
  NAND2_X1 U971 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U972 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U973 ( .A(G160), .B(n867), .ZN(n868) );
  XNOR2_X1 U974 ( .A(n868), .B(n940), .ZN(n885) );
  XNOR2_X1 U975 ( .A(KEYINPUT118), .B(KEYINPUT48), .ZN(n871) );
  XNOR2_X1 U976 ( .A(n869), .B(KEYINPUT46), .ZN(n870) );
  XNOR2_X1 U977 ( .A(n871), .B(n870), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G118), .A2(n527), .ZN(n873) );
  NAND2_X1 U979 ( .A1(G130), .A2(n890), .ZN(n872) );
  NAND2_X1 U980 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n887), .A2(G142), .ZN(n874) );
  XOR2_X1 U982 ( .A(KEYINPUT117), .B(n874), .Z(n876) );
  NAND2_X1 U983 ( .A1(n886), .A2(G106), .ZN(n875) );
  NAND2_X1 U984 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U986 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U987 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U988 ( .A(G164), .B(G162), .ZN(n882) );
  XNOR2_X1 U989 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U990 ( .A(n885), .B(n884), .ZN(n898) );
  NAND2_X1 U991 ( .A1(G103), .A2(n886), .ZN(n889) );
  NAND2_X1 U992 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U993 ( .A1(n889), .A2(n888), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G115), .A2(n527), .ZN(n892) );
  NAND2_X1 U995 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U996 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n952) );
  XNOR2_X1 U999 ( .A(n896), .B(n952), .ZN(n897) );
  XNOR2_X1 U1000 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(G286), .B(G301), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n902), .B(n992), .ZN(n903) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U1006 ( .A(G2454), .B(G2435), .Z(n905) );
  XNOR2_X1 U1007 ( .A(G2438), .B(G2427), .ZN(n904) );
  XNOR2_X1 U1008 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U1009 ( .A(KEYINPUT111), .B(G2446), .Z(n907) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2430), .ZN(n906) );
  XNOR2_X1 U1011 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1012 ( .A(n908), .B(G2451), .Z(n910) );
  XNOR2_X1 U1013 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1014 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1015 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1016 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1025 ( .A(n953), .B(G33), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(n920), .B(G32), .ZN(n921) );
  NAND2_X1 U1027 ( .A1(n922), .A2(n921), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(G25), .B(n923), .ZN(n924) );
  NOR2_X1 U1029 ( .A1(n925), .A2(n924), .ZN(n931) );
  XOR2_X1 U1030 ( .A(G2067), .B(G26), .Z(n926) );
  NAND2_X1 U1031 ( .A1(n926), .A2(G28), .ZN(n929) );
  XOR2_X1 U1032 ( .A(G27), .B(n927), .Z(n928) );
  NOR2_X1 U1033 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1035 ( .A(n932), .B(KEYINPUT53), .ZN(n935) );
  XOR2_X1 U1036 ( .A(G2084), .B(G34), .Z(n933) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NAND2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(G35), .B(G2090), .ZN(n936) );
  NOR2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n965) );
  XNOR2_X1 U1042 ( .A(n938), .B(n965), .ZN(n939) );
  NOR2_X1 U1043 ( .A1(G29), .A2(n939), .ZN(n1024) );
  XNOR2_X1 U1044 ( .A(G160), .B(G2084), .ZN(n941) );
  NAND2_X1 U1045 ( .A1(n941), .A2(n940), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1047 ( .A(KEYINPUT120), .B(n944), .Z(n945) );
  NOR2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n951) );
  INV_X1 U1049 ( .A(n947), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n963) );
  XOR2_X1 U1052 ( .A(G164), .B(G2078), .Z(n955) );
  XNOR2_X1 U1053 ( .A(n953), .B(n952), .ZN(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT50), .B(n956), .ZN(n961) );
  XOR2_X1 U1056 ( .A(G2090), .B(G162), .Z(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1058 ( .A(KEYINPUT51), .B(n959), .Z(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n964), .B(KEYINPUT52), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT122), .B(n967), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n968), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1065 ( .A(G1971), .B(G22), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G23), .B(G1976), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n972) );
  XOR2_X1 U1068 ( .A(G1986), .B(G24), .Z(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n974) );
  XOR2_X1 U1070 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n973) );
  XNOR2_X1 U1071 ( .A(n974), .B(n973), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G21), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G5), .ZN(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(KEYINPUT59), .B(G4), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(n980), .B(n979), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(G20), .B(G1956), .ZN(n981) );
  NOR2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(G1341), .B(G19), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(G1981), .B(G6), .ZN(n983) );
  NOR2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1084 ( .A(KEYINPUT60), .B(n987), .ZN(n988) );
  NOR2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1086 ( .A(KEYINPUT61), .B(n990), .Z(n991) );
  NOR2_X1 U1087 ( .A1(G16), .A2(n991), .ZN(n1019) );
  XNOR2_X1 U1088 ( .A(n992), .B(G1348), .ZN(n1009) );
  XNOR2_X1 U1089 ( .A(G299), .B(G1956), .ZN(n994) );
  XNOR2_X1 U1090 ( .A(G301), .B(G1961), .ZN(n993) );
  NOR2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(G1341), .B(n995), .ZN(n996) );
  NOR2_X1 U1093 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G166), .B(G1971), .ZN(n1000) );
  XOR2_X1 U1096 ( .A(KEYINPUT124), .B(n1000), .Z(n1001) );
  NOR2_X1 U1097 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1099 ( .A(KEYINPUT125), .B(n1005), .Z(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G168), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1104 ( .A(KEYINPUT57), .B(n1012), .Z(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G16), .B(KEYINPUT123), .ZN(n1015) );
  XNOR2_X1 U1107 ( .A(KEYINPUT56), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1020), .Z(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(G11), .ZN(n1026) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

