//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT78), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  OAI211_X1 g010(.A(G128), .B(new_n193), .C1(new_n194), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(new_n199), .C1(KEYINPUT1), .C2(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n214), .A3(KEYINPUT79), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n197), .A2(new_n210), .A3(new_n213), .A4(new_n201), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G134), .ZN(new_n223));
  INV_X1    g037(.A(G134), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n224), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT11), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n222), .A4(G134), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n225), .ZN(new_n232));
  INV_X1    g046(.A(new_n223), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n229), .A2(KEYINPUT65), .A3(new_n230), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n231), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n202), .A2(new_n214), .A3(KEYINPUT10), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT0), .A4(G128), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n198), .A2(new_n199), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n240), .A2(new_n250), .A3(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n242), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n220), .A2(new_n238), .A3(new_n239), .A4(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G110), .B(G140), .ZN(new_n254));
  INV_X1    g068(.A(G227), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G953), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n197), .A2(new_n201), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n210), .A2(new_n213), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n215), .A2(new_n218), .A3(new_n262), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n229), .A2(new_n230), .ZN(new_n264));
  AND4_X1   g078(.A1(KEYINPUT65), .A2(new_n232), .A3(new_n230), .A4(new_n233), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT65), .B1(new_n229), .B2(new_n230), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT81), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n263), .B(new_n267), .C1(new_n268), .C2(KEYINPUT12), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n267), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT12), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n259), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n220), .A2(new_n239), .A3(new_n252), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n267), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n258), .B1(new_n275), .B2(new_n253), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n190), .B(new_n191), .C1(new_n273), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT83), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n253), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n257), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n269), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n253), .A3(new_n258), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n190), .A4(new_n191), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n258), .B1(new_n281), .B2(new_n253), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n275), .A2(new_n253), .A3(new_n258), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT82), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n252), .A2(new_n239), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n216), .B(KEYINPUT79), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n219), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n269), .A2(new_n272), .B1(new_n295), .B2(new_n238), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n292), .B(new_n289), .C1(new_n296), .C2(new_n258), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n190), .B1(new_n298), .B2(new_n191), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n189), .B1(new_n287), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT88), .B(G224), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(G953), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT7), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n260), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n248), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(new_n302), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n246), .B(new_n245), .C1(new_n194), .C2(new_n196), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n304), .B1(new_n309), .B2(new_n243), .ZN(new_n310));
  AOI21_X1  g124(.A(G125), .B1(new_n197), .B2(new_n201), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n303), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(KEYINPUT7), .B(new_n302), .C1(new_n305), .C2(new_n306), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G122), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT8), .Z(new_n316));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G116), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(KEYINPUT5), .ZN(new_n320));
  INV_X1    g134(.A(G116), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G119), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT5), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(new_n318), .A3(KEYINPUT86), .A4(G116), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n320), .A2(new_n323), .A3(G113), .A4(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT2), .B(G113), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G116), .B(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n261), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n214), .A2(new_n330), .A3(new_n326), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n316), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n313), .A2(new_n314), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n331), .A2(new_n261), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n242), .A2(new_n251), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n329), .A2(KEYINPUT66), .A3(KEYINPUT67), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n319), .A2(new_n322), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT66), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n328), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT67), .B1(new_n329), .B2(KEYINPUT66), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n341), .A3(new_n339), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n327), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n336), .B1(new_n337), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT87), .B1(new_n348), .B2(new_n315), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n344), .A2(new_n345), .A3(new_n327), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n327), .B1(new_n344), .B2(new_n345), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n251), .B(new_n242), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(KEYINPUT87), .A3(new_n333), .A4(new_n315), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n335), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(new_n191), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n333), .ZN(new_n357));
  INV_X1    g171(.A(new_n315), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n349), .B2(new_n354), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n308), .A2(new_n312), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n356), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G210), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n352), .A2(new_n333), .A3(new_n315), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT87), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n373), .A2(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n361), .B1(new_n374), .B2(new_n360), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n365), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n356), .A3(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G214), .B1(G237), .B2(G902), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n379), .B(KEYINPUT84), .Z(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT85), .Z(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n300), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G472), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n267), .A2(new_n249), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n224), .A2(G137), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n222), .A2(G134), .ZN(new_n389));
  OAI21_X1  g203(.A(G131), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n197), .A2(new_n201), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n265), .B2(new_n266), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n386), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(new_n386), .C1(new_n238), .C2(new_n248), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n347), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT69), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n350), .A2(new_n351), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT68), .B1(new_n343), .B2(new_n346), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n392), .B1(new_n238), .B2(new_n248), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n236), .A2(new_n237), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n267), .A2(new_n249), .B1(new_n404), .B2(new_n391), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n398), .B1(new_n350), .B2(new_n351), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n343), .A2(KEYINPUT68), .A3(new_n346), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(KEYINPUT69), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(G237), .A2(G953), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G210), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n396), .A2(new_n403), .A3(new_n409), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT31), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n403), .A2(new_n409), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT31), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n414), .A4(new_n396), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT28), .B1(new_n405), .B2(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n402), .A2(new_n347), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n403), .A2(new_n409), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n424), .B2(KEYINPUT28), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(new_n414), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n385), .B(new_n191), .C1(new_n421), .C2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n416), .B(new_n420), .C1(new_n414), .C2(new_n425), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(KEYINPUT32), .A3(new_n385), .A4(new_n191), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n433));
  INV_X1    g247(.A(new_n414), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n402), .A2(KEYINPUT30), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n435), .A2(new_n394), .B1(new_n346), .B2(new_n343), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n417), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n424), .A2(KEYINPUT28), .ZN(new_n438));
  INV_X1    g252(.A(new_n422), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n414), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n433), .B(new_n437), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n403), .B(new_n409), .C1(new_n408), .C2(new_n405), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT28), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n422), .A2(new_n433), .A3(new_n434), .ZN(new_n444));
  AOI21_X1  g258(.A(G902), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT71), .B1(new_n446), .B2(G472), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT71), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n448), .B(new_n385), .C1(new_n441), .C2(new_n445), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n430), .B(new_n432), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n304), .A3(G140), .ZN(new_n452));
  INV_X1    g266(.A(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n304), .A2(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT16), .B(new_n452), .C1(new_n456), .C2(new_n451), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT16), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G146), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT75), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT75), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n463), .A3(G146), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n318), .A2(G128), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n200), .A2(G119), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT72), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT72), .B1(new_n466), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT24), .B(G110), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n466), .B1(KEYINPUT73), .B2(KEYINPUT23), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT23), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n318), .B2(G128), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n478), .A2(G110), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n454), .A2(new_n455), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n195), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n465), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n470), .A2(new_n471), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(G110), .B2(new_n478), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n457), .A2(new_n195), .A3(new_n459), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n461), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G953), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(G221), .A3(G234), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT76), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT22), .B(G137), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n485), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n495), .ZN(new_n497));
  INV_X1    g311(.A(new_n490), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G217), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(G234), .B2(new_n191), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(G902), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n500), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n496), .A2(new_n499), .A3(new_n191), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n505), .B1(new_n511), .B2(new_n502), .ZN(new_n512));
  NAND2_X1  g326(.A1(G234), .A2(G237), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(G952), .A3(new_n491), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(G902), .A3(G953), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT21), .B(G898), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G475), .ZN(new_n520));
  INV_X1    g334(.A(new_n452), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n481), .B2(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G146), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n482), .ZN(new_n524));
  AOI21_X1  g338(.A(G143), .B1(new_n410), .B2(G214), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n410), .A2(G143), .A3(G214), .ZN(new_n527));
  NAND2_X1  g341(.A1(KEYINPUT18), .A2(G131), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n527), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT18), .A3(G131), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n527), .ZN(new_n533));
  OAI21_X1  g347(.A(G131), .B1(new_n533), .B2(new_n525), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n230), .A3(new_n527), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n530), .A2(KEYINPUT17), .A3(G131), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n461), .A2(new_n537), .A3(new_n488), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n532), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G113), .B(G122), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n203), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n532), .A2(new_n539), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n520), .B1(new_n546), .B2(new_n191), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT19), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n456), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n522), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n195), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n534), .A2(new_n535), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n462), .A2(new_n552), .A3(new_n464), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n542), .B1(new_n554), .B2(new_n532), .ZN(new_n555));
  INV_X1    g369(.A(new_n545), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n548), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT20), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT20), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n559), .B(new_n548), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n547), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n188), .A2(new_n501), .A3(G953), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n321), .A2(KEYINPUT14), .A3(G122), .ZN(new_n565));
  XOR2_X1   g379(.A(G116), .B(G122), .Z(new_n566));
  OAI211_X1 g380(.A(G107), .B(new_n565), .C1(new_n566), .C2(KEYINPUT14), .ZN(new_n567));
  XNOR2_X1  g381(.A(G116), .B(G122), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n206), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n200), .A2(G143), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n192), .A2(G128), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n572), .A2(new_n224), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n224), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n567), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n576));
  INV_X1    g390(.A(new_n569), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n568), .A2(new_n206), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n566), .A2(G107), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n569), .A3(KEYINPUT89), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n573), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n571), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n200), .B2(G143), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT90), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n587), .B(new_n583), .C1(new_n200), .C2(G143), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n570), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n584), .B1(new_n589), .B2(KEYINPUT91), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n586), .A2(new_n591), .A3(new_n570), .A4(new_n588), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n224), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n582), .B1(new_n593), .B2(KEYINPUT92), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n570), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n587), .B1(new_n571), .B2(new_n583), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT91), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n584), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G134), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n564), .B(new_n575), .C1(new_n594), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT93), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n593), .A2(KEYINPUT92), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n601), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n582), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT93), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n564), .A4(new_n575), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n575), .B1(new_n594), .B2(new_n602), .ZN(new_n610));
  INV_X1    g424(.A(new_n564), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n604), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT15), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G478), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n191), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n613), .B2(new_n191), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n563), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT94), .A3(new_n616), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n519), .B(new_n562), .C1(new_n619), .C2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n384), .A2(new_n450), .A3(new_n512), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(G101), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G3));
  OAI21_X1  g439(.A(new_n191), .B1(new_n421), .B2(new_n426), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n427), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(KEYINPUT96), .A3(G472), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n512), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n300), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n613), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n610), .B2(new_n611), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n603), .ZN(new_n639));
  INV_X1    g453(.A(G478), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n613), .A2(new_n191), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n640), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n561), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n380), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n355), .A2(new_n191), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n369), .B(new_n647), .C1(new_n375), .C2(new_n365), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n368), .B1(new_n376), .B2(new_n356), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n519), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n378), .A2(KEYINPUT98), .A3(new_n646), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n635), .A2(new_n645), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT99), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n547), .B(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n558), .A2(new_n560), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n619), .A2(new_n664), .A3(new_n621), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n635), .A2(new_n656), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NAND2_X1  g483(.A1(new_n511), .A2(new_n502), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n485), .A2(new_n490), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n503), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n631), .A2(new_n384), .A3(new_n622), .A4(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  AOI21_X1  g492(.A(KEYINPUT98), .B1(new_n378), .B2(new_n646), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n651), .B(new_n380), .C1(new_n370), .C2(new_n377), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n300), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n516), .A2(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n514), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n665), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n685), .A3(new_n450), .A4(new_n675), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  AND3_X1   g501(.A1(new_n619), .A2(new_n621), .A3(new_n562), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n511), .A2(new_n502), .B1(new_n503), .B2(new_n673), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n646), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT105), .Z(new_n691));
  XOR2_X1   g505(.A(new_n683), .B(KEYINPUT39), .Z(new_n692));
  NOR2_X1   g506(.A1(new_n300), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n442), .A2(new_n434), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n415), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n415), .A3(KEYINPUT103), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n191), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT104), .A3(G472), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT104), .B1(new_n702), .B2(G472), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n432), .B(new_n430), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n378), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n691), .A2(new_n695), .A3(new_n696), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  AOI22_X1  g526(.A1(new_n613), .A2(new_n636), .B1(new_n603), .B2(new_n638), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n713), .A2(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n714));
  INV_X1    g528(.A(new_n683), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n714), .A2(KEYINPUT106), .A3(new_n561), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n645), .B2(new_n683), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n681), .A2(new_n450), .A3(new_n675), .A4(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT107), .B(G146), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G48));
  NOR2_X1   g536(.A1(new_n679), .A2(new_n680), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n653), .A3(new_n645), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n283), .A2(new_n191), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n286), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n189), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n450), .A2(new_n512), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT41), .B(G113), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND4_X1  g547(.A1(new_n665), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n321), .ZN(G18));
  NAND3_X1  g550(.A1(new_n450), .A2(new_n622), .A3(new_n675), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n652), .A2(new_n729), .A3(new_n654), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n318), .ZN(G21));
  AND2_X1   g554(.A1(new_n416), .A2(new_n420), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n422), .B1(new_n442), .B2(KEYINPUT28), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n434), .B1(new_n742), .B2(KEYINPUT108), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(G472), .A2(G902), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n746), .A2(new_n747), .B1(new_n626), .B2(G472), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n688), .A3(new_n729), .A4(new_n512), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n655), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(G122), .Z(G24));
  INV_X1    g565(.A(new_n738), .ZN(new_n752));
  INV_X1    g566(.A(new_n747), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n443), .A2(new_n439), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n434), .A3(new_n743), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n757), .B2(new_n741), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n385), .B1(new_n431), .B2(new_n191), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n689), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n752), .A2(new_n719), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n289), .B1(new_n296), .B2(new_n258), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n190), .B1(new_n765), .B2(new_n191), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n728), .B1(new_n286), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n370), .A2(new_n377), .A3(new_n646), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n370), .A2(new_n377), .A3(new_n646), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n768), .A3(KEYINPUT109), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n763), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT32), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n427), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n776), .B(new_n432), .C1(new_n447), .C2(new_n449), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n512), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT110), .B1(new_n777), .B2(new_n512), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n719), .B(new_n774), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n766), .B1(new_n278), .B2(new_n285), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n770), .A2(new_n781), .A3(new_n764), .A4(new_n728), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT109), .B1(new_n772), .B2(new_n768), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n450), .B(new_n512), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n719), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n763), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  OR2_X1    g602(.A1(new_n784), .A2(new_n684), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  NAND2_X1  g604(.A1(new_n642), .A2(new_n644), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n561), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT43), .Z(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n630), .A3(new_n629), .A4(new_n675), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT111), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n291), .B2(new_n297), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n799));
  OAI21_X1  g613(.A(G469), .B1(new_n765), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(G469), .A2(G902), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT46), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n287), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n189), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n692), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n794), .A2(new_n795), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n772), .B(KEYINPUT112), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n797), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(KEYINPUT47), .A3(new_n189), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n450), .A2(new_n512), .A3(new_n770), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n719), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT113), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND2_X1  g635(.A1(new_n748), .A2(new_n512), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n793), .A2(new_n515), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n793), .A2(new_n825), .A3(new_n515), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n709), .A2(new_n380), .A3(new_n729), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n727), .A2(new_n189), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n811), .B(new_n827), .C1(new_n817), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n729), .A2(new_n772), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n632), .A3(new_n514), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n707), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n562), .A3(new_n791), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n834), .B1(new_n824), .B2(new_n826), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n760), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n831), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT51), .ZN(new_n841));
  INV_X1    g655(.A(new_n645), .ZN(new_n842));
  OAI211_X1 g656(.A(G952), .B(new_n491), .C1(new_n836), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n752), .B2(new_n827), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n778), .A2(new_n779), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n846), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT119), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n686), .A2(new_n761), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n769), .A2(new_n675), .A3(new_n715), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n706), .A2(new_n856), .A3(new_n723), .A4(new_n688), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n720), .A2(new_n857), .A3(KEYINPUT52), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n686), .A2(new_n761), .A3(KEYINPUT115), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n686), .A2(new_n720), .A3(new_n761), .A4(new_n857), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n719), .B(new_n760), .C1(new_n783), .C2(new_n782), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n617), .A2(new_n618), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n664), .A2(new_n868), .A3(new_n683), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n300), .A2(new_n869), .A3(new_n770), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n450), .A3(new_n675), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n867), .B(new_n871), .C1(new_n784), .C2(new_n684), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n786), .B2(new_n780), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n842), .B1(new_n868), .B2(new_n562), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n383), .A2(new_n519), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n631), .A2(new_n633), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n676), .A2(new_n876), .A3(new_n623), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n730), .B1(new_n724), .B2(new_n734), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n737), .A2(new_n738), .B1(new_n655), .B2(new_n749), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n873), .A2(new_n880), .ZN(new_n885));
  INV_X1    g699(.A(new_n853), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n858), .A2(new_n886), .B1(new_n861), .B2(new_n863), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n882), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n885), .A2(new_n887), .A3(new_n884), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT114), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n873), .A2(new_n880), .A3(KEYINPUT114), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n866), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n895), .B2(new_n883), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n852), .A2(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n709), .A2(new_n512), .A3(new_n189), .A4(new_n382), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n727), .B(KEYINPUT49), .ZN(new_n899));
  OR4_X1    g713(.A1(new_n706), .A2(new_n898), .A3(new_n792), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n491), .A2(G952), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT121), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n873), .A2(new_n880), .A3(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n861), .A2(new_n863), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT116), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n860), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n858), .A2(new_n886), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n906), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT53), .B1(new_n881), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n191), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n375), .B(new_n366), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n919), .B(new_n920), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n916), .A2(new_n917), .A3(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n904), .B1(new_n923), .B2(new_n924), .ZN(G51));
  AOI21_X1  g739(.A(KEYINPUT123), .B1(new_n915), .B2(new_n801), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n914), .A2(new_n927), .A3(new_n191), .A4(new_n802), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT54), .B1(new_n910), .B2(new_n913), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n889), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n803), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n283), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n902), .B1(new_n929), .B2(new_n935), .ZN(G54));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n937));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n915), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n555), .A2(new_n556), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n902), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  INV_X1    g756(.A(new_n940), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n915), .A2(KEYINPUT124), .A3(new_n943), .A4(new_n938), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(G60));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n713), .B1(new_n896), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n713), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n910), .A2(new_n913), .A3(KEYINPUT54), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n883), .B1(new_n882), .B2(new_n888), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n903), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n946), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n904), .B1(new_n931), .B2(new_n951), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n873), .A2(KEYINPUT114), .A3(new_n880), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT114), .B1(new_n873), .B2(new_n880), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n960), .B2(new_n866), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT54), .B1(new_n961), .B2(new_n890), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n948), .B1(new_n962), .B2(new_n889), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT125), .B(new_n957), .C1(new_n963), .C2(new_n713), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n956), .A2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n914), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n673), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n500), .B1(new_n914), .B2(new_n967), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n903), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n969), .A2(KEYINPUT61), .A3(new_n903), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G66));
  OAI21_X1  g789(.A(G953), .B1(new_n518), .B2(new_n301), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n880), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n364), .B1(G898), .B2(new_n491), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  NOR2_X1   g793(.A1(new_n393), .A2(new_n395), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n551), .B(KEYINPUT126), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n855), .A2(new_n720), .A3(new_n859), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n820), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n809), .A2(new_n845), .A3(new_n723), .A4(new_n688), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n812), .A2(new_n985), .A3(new_n787), .A4(new_n789), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n491), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n255), .A2(G900), .A3(G953), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n694), .A2(new_n770), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n874), .B(KEYINPUT127), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n991), .A2(new_n992), .A3(new_n450), .A4(new_n512), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n820), .A2(new_n812), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n983), .A2(new_n711), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n990), .B1(new_n998), .B2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n989), .B1(new_n999), .B2(new_n982), .ZN(G72));
  NOR3_X1   g814(.A1(new_n417), .A2(new_n436), .A3(new_n414), .ZN(new_n1001));
  INV_X1    g815(.A(new_n880), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n984), .A2(new_n986), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n902), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n414), .B1(new_n417), .B2(new_n436), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n994), .A2(new_n880), .A3(new_n996), .A4(new_n997), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n1005), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1006), .B(new_n895), .C1(new_n437), .C2(new_n415), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(G57));
endmodule


