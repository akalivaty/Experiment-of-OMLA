//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G99gat), .ZN(new_n205));
  INV_X1    g004(.A(G106gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT8), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT97), .B(G92gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G85gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT98), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT7), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G99gat), .B(G106gat), .Z(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G57gat), .B(G64gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT92), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT93), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G71gat), .B(G78gat), .Z(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT91), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n217), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n221), .A2(new_n223), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n215), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(KEYINPUT101), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT10), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n216), .A2(new_n227), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n216), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(KEYINPUT10), .A3(new_n225), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n204), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n204), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(new_n228), .B2(new_n230), .ZN(new_n236));
  XNOR2_X1  g035(.A(G120gat), .B(G148gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G176gat), .B(G204gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  OR3_X1    g038(.A1(new_n234), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n234), .B2(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n225), .A2(KEYINPUT21), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT94), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n245));
  XNOR2_X1  g044(.A(G183gat), .B(G211gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n244), .B(new_n247), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n225), .A2(KEYINPUT21), .ZN(new_n250));
  XOR2_X1   g049(.A(G15gat), .B(G22gat), .Z(new_n251));
  INV_X1    g050(.A(G1gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(G8gat), .B1(new_n253), .B2(KEYINPUT89), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n252), .A2(KEYINPUT16), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n255), .B2(new_n251), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n254), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT95), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G155gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(G155gat), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G231gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(new_n203), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n267), .A2(new_n270), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n249), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n273), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n271), .A3(new_n248), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT15), .ZN(new_n277));
  XOR2_X1   g076(.A(G43gat), .B(G50gat), .Z(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT88), .ZN(new_n279));
  NAND2_X1  g078(.A1(G29gat), .A2(G36gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT14), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G29gat), .B2(G36gat), .ZN(new_n282));
  INV_X1    g081(.A(G29gat), .ZN(new_n283));
  INV_X1    g082(.A(G36gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT14), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n280), .A3(new_n282), .A4(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n282), .A3(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n278), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n277), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(KEYINPUT88), .B2(new_n278), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT15), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n232), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(KEYINPUT17), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n216), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G190gat), .B(G218gat), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT99), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n297), .B(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(G162gat), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT96), .B(G134gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT100), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n297), .A2(new_n299), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n307), .B2(KEYINPUT100), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n300), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n274), .A2(new_n276), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n313));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT4), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n317), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n318), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT71), .B(KEYINPUT2), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n325), .B(new_n326), .C1(new_n317), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(KEYINPUT71), .A2(KEYINPUT2), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT71), .A2(KEYINPUT2), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(G148gat), .ZN(new_n333));
  INV_X1    g132(.A(G148gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(G141gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n330), .B(new_n331), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n326), .B1(new_n336), .B2(new_n325), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n323), .B1(new_n329), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G120gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G113gat), .ZN(new_n340));
  INV_X1    g139(.A(G113gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G120gat), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT1), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT65), .B(G134gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT66), .B(G127gat), .ZN(new_n348));
  INV_X1    g147(.A(G134gat), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n260), .A2(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT4), .B1(new_n338), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n325), .B1(new_n317), .B2(new_n327), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT72), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n322), .B1(new_n356), .B2(new_n328), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n338), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n323), .B(new_n367), .C1(new_n329), .C2(new_n337), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n353), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n316), .B(new_n361), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n359), .B1(new_n364), .B2(new_n365), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n338), .A2(new_n353), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n315), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(KEYINPUT5), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n361), .B(new_n375), .C1(new_n366), .C2(new_n369), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  INV_X1    g183(.A(new_n382), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n374), .A2(new_n385), .A3(new_n376), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n374), .B2(new_n376), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT6), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  XNOR2_X1  g190(.A(G197gat), .B(G204gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT22), .ZN(new_n393));
  INV_X1    g192(.A(G211gat), .ZN(new_n394));
  INV_X1    g193(.A(G218gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G211gat), .B(G218gat), .Z(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  NOR2_X1   g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT23), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G169gat), .ZN(new_n405));
  INV_X1    g204(.A(G176gat), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT23), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G183gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT64), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G183gat), .ZN(new_n412));
  AOI21_X1  g211(.A(G190gat), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT24), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n404), .B(new_n408), .C1(new_n413), .C2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT25), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n407), .B1(new_n401), .B2(new_n403), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n419), .A2(KEYINPUT25), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n410), .A2(new_n412), .A3(KEYINPUT27), .ZN(new_n429));
  NOR2_X1   g228(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(KEYINPUT27), .B(G183gat), .Z(new_n432));
  OAI21_X1  g231(.A(KEYINPUT28), .B1(new_n432), .B2(G190gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT26), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n400), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n402), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n431), .A2(new_n433), .A3(new_n414), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n427), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n427), .B2(new_n438), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n399), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n443), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n397), .B(new_n398), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n445), .B(new_n446), .C1(new_n441), .C2(new_n439), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G8gat), .B(G36gat), .ZN(new_n449));
  INV_X1    g248(.A(G92gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT70), .B(G64gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n391), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n454), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n444), .A2(KEYINPUT30), .A3(new_n447), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT76), .B1(new_n390), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n461), .B(new_n458), .C1(new_n387), .C2(new_n389), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT29), .B1(new_n357), .B2(new_n367), .ZN(new_n463));
  INV_X1    g262(.A(new_n367), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n446), .B2(new_n465), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n463), .A2(new_n446), .B1(new_n357), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT78), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n368), .A2(new_n470), .A3(new_n465), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n368), .B2(new_n465), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(new_n446), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n362), .B1(new_n399), .B2(KEYINPUT29), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n363), .B(new_n322), .C1(new_n356), .C2(new_n328), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n468), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n469), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT79), .B1(new_n480), .B2(G22gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G78gat), .B(G106gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G50gat), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT77), .B(KEYINPUT31), .Z(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n480), .A2(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(G22gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n463), .A2(new_n470), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n368), .A2(new_n465), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT78), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(new_n399), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n478), .A3(new_n477), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n488), .B1(new_n493), .B2(new_n469), .ZN(new_n494));
  OAI22_X1  g293(.A1(new_n481), .A2(new_n486), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n480), .A2(G22gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n488), .A3(new_n469), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT79), .A4(new_n485), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n427), .A2(new_n359), .A3(new_n438), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n427), .A2(new_n438), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n353), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n427), .A2(new_n359), .A3(new_n438), .A4(KEYINPUT67), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G43gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G71gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n205), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n509), .B(KEYINPUT32), .C1(new_n511), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n502), .A2(new_n507), .A3(new_n504), .A4(new_n505), .ZN(new_n520));
  OR3_X1    g319(.A1(new_n520), .A2(KEYINPUT68), .A3(KEYINPUT34), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT68), .B1(new_n520), .B2(KEYINPUT34), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n519), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n519), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n499), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n460), .A2(new_n462), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n313), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT82), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n387), .A2(new_n532), .B1(KEYINPUT85), .B2(new_n389), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n389), .A2(KEYINPUT85), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n374), .A2(new_n385), .A3(new_n376), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n535), .A2(new_n388), .A3(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT82), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n499), .ZN(new_n539));
  INV_X1    g338(.A(new_n524), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n519), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n518), .A3(new_n516), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n458), .B(KEYINPUT80), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n538), .A2(new_n544), .A3(new_n530), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n389), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n459), .B1(new_n536), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n461), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n390), .A2(KEYINPUT76), .A3(new_n459), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n519), .A2(new_n525), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n540), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n519), .A2(new_n524), .A3(new_n525), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(new_n498), .B2(new_n495), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n531), .A2(new_n547), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n361), .B1(new_n366), .B2(new_n369), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n561), .B2(new_n314), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(KEYINPUT81), .A3(new_n315), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT39), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n371), .A2(new_n372), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n565), .B1(new_n567), .B2(new_n314), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n385), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n566), .A2(KEYINPUT40), .A3(new_n385), .A4(new_n569), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n545), .A3(new_n383), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n447), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT37), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n447), .A4(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(new_n577), .A3(new_n454), .A4(new_n579), .ZN(new_n580));
  OAI22_X1  g379(.A1(new_n580), .A2(KEYINPUT84), .B1(new_n454), .B2(new_n448), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(KEYINPUT84), .B2(new_n580), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n534), .A3(new_n533), .A4(new_n537), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n576), .A2(new_n579), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n577), .B1(new_n584), .B2(new_n454), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n574), .B(new_n499), .C1(new_n583), .C2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n539), .B1(new_n460), .B2(new_n462), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n526), .A2(new_n527), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n543), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AOI211_X1 g391(.A(new_n242), .B(new_n312), .C1(new_n558), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n294), .A2(new_n257), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR3_X1    g395(.A1(new_n257), .A2(new_n289), .A3(new_n291), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n294), .A2(KEYINPUT90), .A3(new_n257), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT18), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n292), .B(new_n257), .Z(new_n602));
  XOR2_X1   g401(.A(new_n598), .B(KEYINPUT13), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  INV_X1    g405(.A(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT11), .B(G169gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT87), .Z(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT12), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n601), .A2(new_n612), .A3(new_n604), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n593), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n390), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n252), .ZN(G1324gat));
  INV_X1    g418(.A(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n545), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT42), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT16), .B(G8gat), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT103), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n621), .B(KEYINPUT102), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n622), .B1(new_n626), .B2(G8gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n623), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(G1325gat));
  INV_X1    g428(.A(G15gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n591), .B(KEYINPUT104), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n617), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n620), .A2(new_n590), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n630), .B2(new_n633), .ZN(G1326gat));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n499), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT43), .B(G22gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1327gat));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n311), .A2(KEYINPUT44), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n558), .A2(KEYINPUT106), .A3(new_n592), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT106), .B1(new_n558), .B2(new_n592), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n556), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT86), .B1(new_n556), .B2(KEYINPUT35), .ZN(new_n644));
  INV_X1    g443(.A(new_n547), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n310), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651));
  INV_X1    g450(.A(new_n615), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n612), .B1(new_n601), .B2(new_n604), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n614), .A2(KEYINPUT105), .A3(new_n615), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n274), .A2(new_n276), .ZN(new_n658));
  INV_X1    g457(.A(new_n242), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n638), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  AOI211_X1 g461(.A(KEYINPUT107), .B(new_n660), .C1(new_n642), .C2(new_n649), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664), .B2(new_n390), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n652), .A2(new_n653), .ZN(new_n666));
  INV_X1    g465(.A(new_n658), .ZN(new_n667));
  NOR4_X1   g466(.A1(new_n648), .A2(new_n666), .A3(new_n667), .A4(new_n242), .ZN(new_n668));
  INV_X1    g467(.A(new_n390), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n283), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(new_n671), .ZN(G1328gat));
  OAI21_X1  g471(.A(G36gat), .B1(new_n664), .B2(new_n546), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n284), .A3(new_n545), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(KEYINPUT46), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(KEYINPUT108), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT46), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n678), .A3(new_n679), .ZN(G1329gat));
  INV_X1    g479(.A(G43gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n668), .A2(new_n681), .A3(new_n590), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n631), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n662), .B2(new_n663), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(G43gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n639), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n646), .B2(new_n647), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n558), .A2(KEYINPUT106), .A3(new_n592), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n311), .B1(new_n558), .B2(new_n592), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n661), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G43gat), .B1(new_n696), .B2(new_n591), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n683), .B1(new_n697), .B2(new_n682), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n687), .A2(KEYINPUT109), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  INV_X1    g499(.A(new_n684), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n650), .A2(new_n638), .A3(new_n661), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n631), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(new_n681), .ZN(new_n705));
  INV_X1    g504(.A(new_n698), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n699), .A2(new_n707), .ZN(G1330gat));
  OAI21_X1  g507(.A(G50gat), .B1(new_n696), .B2(new_n499), .ZN(new_n709));
  INV_X1    g508(.A(G50gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n668), .A2(new_n710), .A3(new_n539), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(KEYINPUT48), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n711), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n539), .B1(new_n662), .B2(new_n663), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(G50gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n715), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n312), .A2(new_n657), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n242), .B(new_n717), .C1(new_n640), .C2(new_n641), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n669), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n546), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(G1333gat));
  OR3_X1    g529(.A1(new_n722), .A2(G71gat), .A3(new_n543), .ZN(new_n731));
  OAI21_X1  g530(.A(G71gat), .B1(new_n722), .B2(new_n631), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n539), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  XNOR2_X1  g537(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n739));
  NAND2_X1  g538(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n667), .A2(new_n657), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n693), .A2(new_n741), .ZN(new_n742));
  MUX2_X1   g541(.A(new_n739), .B(new_n740), .S(new_n742), .Z(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n242), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n669), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n650), .A2(new_n242), .A3(new_n741), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n669), .A2(G85gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  INV_X1    g548(.A(new_n208), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n545), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n742), .A2(KEYINPUT112), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n545), .A2(new_n450), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n659), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n744), .B2(new_n754), .ZN(new_n758));
  OAI22_X1  g557(.A1(new_n756), .A2(new_n757), .B1(new_n751), .B2(new_n758), .ZN(G1337gat));
  INV_X1    g558(.A(new_n747), .ZN(new_n760));
  OAI21_X1  g559(.A(G99gat), .B1(new_n760), .B2(new_n631), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n590), .A2(new_n205), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n744), .B2(new_n762), .ZN(G1338gat));
  OAI21_X1  g562(.A(G106gat), .B1(new_n760), .B2(new_n499), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n659), .A2(G106gat), .A3(new_n499), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT53), .B1(new_n743), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n753), .A2(new_n765), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  NAND2_X1  g570(.A1(new_n717), .A2(new_n659), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n773), .A2(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n610), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n310), .A2(new_n615), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n231), .A2(new_n233), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n235), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n239), .B1(new_n779), .B2(KEYINPUT54), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n231), .A2(new_n204), .A3(new_n233), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT54), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n234), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n239), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n234), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(KEYINPUT55), .C1(new_n234), .C2(new_n782), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n240), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n784), .A2(KEYINPUT113), .A3(new_n240), .A4(new_n788), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n776), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n615), .A2(new_n242), .A3(new_n775), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n656), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n793), .B1(new_n796), .B2(new_n311), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n772), .B1(new_n797), .B2(new_n667), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n545), .A2(new_n390), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n798), .A2(new_n555), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n341), .A3(new_n657), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n544), .A3(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n666), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1340gat));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n339), .A3(new_n242), .ZN(new_n805));
  OAI21_X1  g604(.A(G120gat), .B1(new_n802), .B2(new_n659), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1341gat));
  AOI21_X1  g606(.A(new_n348), .B1(new_n800), .B2(new_n667), .ZN(new_n808));
  INV_X1    g607(.A(new_n348), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n802), .A2(new_n809), .A3(new_n658), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(G1342gat));
  INV_X1    g610(.A(new_n347), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n800), .A2(new_n812), .A3(new_n310), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT56), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n813), .A2(KEYINPUT56), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n802), .B2(new_n311), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(G1343gat));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n539), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n685), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n666), .A2(G141gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT116), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(new_n799), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(KEYINPUT117), .B2(KEYINPUT58), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n615), .A2(new_n242), .A3(new_n775), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n784), .A2(new_n240), .A3(new_n788), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n616), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(new_n310), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n776), .A2(new_n791), .A3(new_n792), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n794), .B1(new_n666), .B2(new_n789), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n311), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n835), .A2(new_n658), .B1(new_n659), .B2(new_n717), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT57), .B1(new_n836), .B2(new_n499), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n798), .A2(new_n838), .A3(new_n539), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n591), .A2(new_n799), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n826), .B1(new_n841), .B2(new_n666), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n825), .B1(new_n332), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n841), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n332), .B1(new_n844), .B2(new_n657), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(KEYINPUT117), .B2(new_n824), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n826), .ZN(G1344gat));
  NAND4_X1  g646(.A1(new_n821), .A2(new_n334), .A3(new_n242), .A4(new_n799), .ZN(new_n848));
  XOR2_X1   g647(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n849));
  NAND2_X1  g648(.A1(new_n820), .A2(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n311), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n776), .A2(new_n829), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n667), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n312), .A2(new_n616), .A3(new_n242), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n838), .B(new_n539), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n850), .A2(new_n242), .A3(new_n840), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n849), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n837), .A2(new_n839), .A3(new_n242), .A4(new_n840), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n858), .A2(new_n859), .A3(G148gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n848), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT119), .B(new_n848), .C1(new_n857), .C2(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1345gat));
  NOR3_X1   g664(.A1(new_n841), .A2(new_n264), .A3(new_n658), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n821), .A2(new_n667), .A3(new_n799), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n264), .B2(new_n867), .ZN(G1346gat));
  NAND3_X1  g667(.A1(new_n844), .A2(G162gat), .A3(new_n310), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n821), .A2(new_n310), .A3(new_n799), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(G162gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n869), .B(KEYINPUT120), .C1(new_n870), .C2(G162gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n546), .A2(new_n669), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n798), .A2(new_n555), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n405), .A3(new_n657), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT121), .Z(new_n879));
  NAND3_X1  g678(.A1(new_n798), .A2(new_n544), .A3(new_n876), .ZN(new_n880));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n666), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT122), .Z(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(G1348gat));
  AOI21_X1  g682(.A(G176gat), .B1(new_n877), .B2(new_n242), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n880), .A2(new_n406), .A3(new_n659), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(G1349gat));
  INV_X1    g685(.A(new_n432), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n877), .A2(new_n667), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n410), .B(new_n412), .C1(new_n880), .C2(new_n658), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n880), .B2(new_n311), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n423), .A3(new_n310), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1351gat));
  AND2_X1   g696(.A1(new_n821), .A2(new_n876), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n607), .A3(new_n657), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n631), .A2(new_n876), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n850), .A2(new_n855), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G197gat), .B1(new_n902), .B2(new_n666), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n903), .ZN(G1352gat));
  NAND3_X1  g703(.A1(new_n821), .A2(new_n242), .A3(new_n876), .ZN(new_n905));
  XOR2_X1   g704(.A(KEYINPUT125), .B(G204gat), .Z(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT62), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n850), .A2(new_n855), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n242), .A3(new_n901), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT126), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n909), .A2(new_n912), .A3(new_n242), .A4(new_n901), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n908), .A2(new_n914), .ZN(G1353gat));
  OAI21_X1  g714(.A(G211gat), .B1(new_n902), .B2(new_n658), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT63), .B(G211gat), .C1(new_n902), .C2(new_n658), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(KEYINPUT127), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n394), .A3(new_n667), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n916), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(G1354gat));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n395), .A3(new_n310), .ZN(new_n925));
  OAI21_X1  g724(.A(G218gat), .B1(new_n902), .B2(new_n311), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


