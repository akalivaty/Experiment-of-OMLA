//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G211gat), .B2(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n202), .B2(new_n203), .ZN(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n205), .B2(new_n207), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211));
  NAND2_X1  g010(.A1(G226gat), .A2(G233gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT27), .B(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT28), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT27), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT27), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G183gat), .ZN(new_n230));
  AND4_X1   g029(.A1(KEYINPUT28), .A2(new_n228), .A3(new_n230), .A4(new_n225), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n223), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(G190gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n216), .B1(KEYINPUT23), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(KEYINPUT23), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(KEYINPUT25), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n221), .A2(new_n245), .A3(new_n236), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n221), .B2(new_n236), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n235), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n235), .B(new_n250), .C1(new_n246), .C2(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n240), .A2(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n218), .A2(new_n219), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n215), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n241), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n249), .A2(new_n251), .A3(new_n252), .A4(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n244), .B1(KEYINPUT25), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n212), .B1(new_n259), .B2(KEYINPUT29), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(KEYINPUT25), .ZN(new_n261));
  INV_X1    g060(.A(new_n244), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n212), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n211), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT72), .B1(new_n263), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n210), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n260), .A2(new_n265), .ZN(new_n269));
  INV_X1    g068(.A(new_n210), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT73), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279));
  AOI211_X1 g078(.A(new_n279), .B(new_n275), .C1(new_n268), .C2(new_n271), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n268), .A2(new_n271), .A3(new_n275), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(KEYINPUT30), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n278), .A2(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G127gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G134gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G127gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT67), .ZN(new_n290));
  OR3_X1    g089(.A1(new_n288), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G113gat), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G120gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT1), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n294), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n300), .A2(new_n287), .A3(new_n289), .A4(new_n301), .ZN(new_n302));
  OAI22_X1  g101(.A1(new_n292), .A2(new_n297), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n263), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G227gat), .A2(G233gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n259), .A2(new_n303), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G71gat), .B(G99gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT69), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n312), .B(G15gat), .Z(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(G43gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT34), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI211_X1 g118(.A(KEYINPUT34), .B(new_n306), .C1(new_n305), .C2(new_n307), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n308), .A2(KEYINPUT32), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n317), .A2(new_n318), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n310), .B(new_n315), .C1(new_n324), .C2(new_n320), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n323), .B1(new_n322), .B2(new_n325), .ZN(new_n327));
  XOR2_X1   g126(.A(G78gat), .B(G106gat), .Z(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G50gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G141gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT74), .B(G141gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(KEYINPUT2), .ZN(new_n343));
  XNOR2_X1  g142(.A(G155gat), .B(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n336), .A2(new_n342), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  XNOR2_X1  g146(.A(G141gat), .B(G148gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n341), .B(new_n339), .C1(new_n348), .C2(KEYINPUT2), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n270), .B1(new_n332), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n342), .A3(new_n343), .ZN(new_n352));
  INV_X1    g151(.A(new_n334), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT74), .B(G141gat), .Z(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(G148gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n332), .B1(new_n208), .B2(new_n209), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  INV_X1    g158(.A(G228gat), .ZN(new_n360));
  INV_X1    g159(.A(G233gat), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n351), .A2(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n350), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n210), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n360), .A2(new_n361), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n358), .A2(new_n347), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n365), .C1(new_n357), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT84), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G22gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n331), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n370), .A3(G22gat), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT83), .B(G22gat), .Z(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n331), .ZN(new_n376));
  NOR2_X1   g175(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n368), .B2(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n372), .A2(new_n373), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n326), .A2(new_n327), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT6), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n303), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n294), .A2(new_n296), .A3(new_n298), .ZN(new_n390));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n390), .A2(new_n301), .A3(new_n391), .A4(new_n300), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n392), .B(KEYINPUT76), .C1(new_n297), .C2(new_n292), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n387), .A2(new_n350), .A3(new_n389), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT4), .B1(new_n356), .B2(new_n303), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n304), .A2(new_n399), .A3(new_n346), .A4(new_n349), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n357), .A2(new_n304), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT77), .ZN(new_n407));
  AND4_X1   g206(.A1(new_n395), .A2(new_n406), .A3(new_n407), .A4(new_n394), .ZN(new_n408));
  INV_X1    g207(.A(new_n395), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n356), .A3(new_n393), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n389), .A2(new_n356), .A3(KEYINPUT78), .A4(new_n393), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n409), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n397), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n411), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n404), .A3(new_n413), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n397), .B1(new_n421), .B2(new_n409), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT80), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n403), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n407), .A3(new_n406), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n422), .B2(KEYINPUT80), .ZN(new_n426));
  AOI211_X1 g225(.A(new_n418), .B(new_n397), .C1(new_n421), .C2(new_n409), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n426), .A2(KEYINPUT81), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n402), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n384), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n386), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n402), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT81), .B1(new_n426), .B2(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n418), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n437), .A2(new_n403), .A3(new_n423), .A4(new_n425), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n439), .A2(new_n432), .A3(new_n385), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n285), .B(new_n380), .C1(new_n434), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n442), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n282), .A2(KEYINPUT30), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n282), .A2(KEYINPUT30), .ZN(new_n447));
  OAI22_X1  g246(.A1(new_n446), .A2(new_n447), .B1(new_n277), .B2(new_n280), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n386), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(new_n431), .A3(new_n430), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(KEYINPUT86), .A3(new_n380), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(KEYINPUT35), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n395), .B1(new_n401), .B2(new_n394), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n409), .B2(new_n421), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n430), .B1(new_n454), .B2(new_n455), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT40), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n448), .B(new_n460), .C1(new_n439), .C2(new_n384), .ZN(new_n461));
  INV_X1    g260(.A(new_n379), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n272), .A2(new_n276), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n276), .A2(KEYINPUT37), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n272), .A2(KEYINPUT37), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT38), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n282), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n269), .B2(new_n210), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n270), .B1(new_n266), .B2(new_n267), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT38), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n466), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n450), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n470), .B1(new_n477), .B2(KEYINPUT85), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n449), .A2(new_n476), .A3(new_n479), .A4(new_n450), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n463), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT36), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n326), .A2(new_n327), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT70), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT70), .B(KEYINPUT36), .C1(new_n326), .C2(new_n327), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n485), .B(new_n486), .C1(new_n451), .C2(new_n462), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n444), .B(new_n453), .C1(new_n481), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G36gat), .ZN(new_n489));
  AND2_X1   g288(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G29gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n497));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT17), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(G1gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  OR2_X1    g303(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n503), .B2(KEYINPUT90), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n512), .A2(new_n514), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT91), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT91), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n500), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n522), .ZN(new_n523));
  OR3_X1    g322(.A1(new_n500), .A2(new_n515), .A3(new_n516), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n520), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n522), .B(KEYINPUT13), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(new_n522), .A3(new_n520), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n523), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G169gat), .B(G197gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT12), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n527), .A3(new_n530), .A4(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n488), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n449), .A2(new_n450), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G57gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G64gat), .ZN(new_n546));
  INV_X1    g345(.A(G64gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(KEYINPUT9), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(G71gat), .A2(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n555), .A3(new_n550), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g356(.A(new_n553), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n550), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT93), .B1(new_n551), .B2(new_n553), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n557), .A2(new_n560), .A3(new_n561), .A4(new_n549), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n286), .ZN(new_n568));
  INV_X1    g367(.A(new_n563), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n516), .B(new_n515), .C1(KEYINPUT21), .C2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n337), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n586));
  XNOR2_X1  g385(.A(G99gat), .B(G106gat), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n581), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n586), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n569), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n588), .B(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n563), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n597), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n591), .A2(new_n594), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G230gat), .A3(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G120gat), .B(G148gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT97), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n608), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n501), .A2(new_n593), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n590), .A2(new_n500), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n613), .B2(new_n615), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G134gat), .B(G162gat), .Z(new_n622));
  NOR2_X1   g421(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n624), .B(KEYINPUT95), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n619), .B2(new_n620), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n579), .A2(new_n612), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n542), .A2(new_n544), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n285), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n513), .B1(new_n542), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT98), .Z(new_n637));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n542), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT42), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(G1325gat));
  NAND2_X1  g440(.A1(new_n542), .A2(new_n632), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(G15gat), .B1(new_n643), .B2(new_n483), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n485), .A2(new_n486), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G15gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT99), .Z(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n643), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n642), .A2(new_n462), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT43), .B(G22gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  INV_X1    g450(.A(new_n612), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(new_n579), .A3(new_n630), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n542), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n493), .A3(new_n544), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT45), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n579), .B(KEYINPUT100), .Z(new_n658));
  AND3_X1   g457(.A1(new_n658), .A2(new_n541), .A3(new_n612), .ZN(new_n659));
  INV_X1    g458(.A(new_n630), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT44), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n453), .A2(new_n444), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n477), .A2(KEYINPUT85), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n480), .A3(new_n469), .ZN(new_n665));
  INV_X1    g464(.A(new_n463), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n487), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n660), .B(new_n662), .C1(new_n663), .C2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n488), .B2(new_n660), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n659), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n674), .B(new_n659), .C1(new_n669), .C2(new_n671), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n673), .A2(new_n544), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n657), .B1(new_n493), .B2(new_n676), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n655), .A2(new_n489), .A3(new_n448), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n673), .A2(new_n448), .A3(new_n675), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G36gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(new_n483), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n654), .A2(G43gat), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n645), .ZN(new_n689));
  OAI21_X1  g488(.A(G43gat), .B1(new_n672), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(KEYINPUT47), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n645), .A3(new_n675), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n692), .A2(new_n693), .A3(G43gat), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n692), .B2(G43gat), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n694), .A2(new_n695), .A3(new_n687), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n691), .B1(new_n696), .B2(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g496(.A1(new_n672), .A2(KEYINPUT105), .A3(new_n462), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT105), .B1(new_n672), .B2(new_n462), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(G50gat), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n654), .A2(G50gat), .A3(new_n462), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(KEYINPUT48), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n700), .B2(new_n703), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n673), .A2(new_n379), .A3(new_n675), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G50gat), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(new_n702), .ZN(new_n708));
  OAI22_X1  g507(.A1(new_n704), .A2(new_n705), .B1(new_n708), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g508(.A(new_n541), .ZN(new_n710));
  INV_X1    g509(.A(new_n579), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n660), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n710), .A2(new_n488), .A3(new_n712), .A4(new_n652), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n543), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n545), .ZN(G1332gat));
  NOR2_X1   g517(.A1(new_n716), .A2(new_n285), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  AND2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n719), .B2(new_n720), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n716), .B2(new_n689), .ZN(new_n724));
  INV_X1    g523(.A(G71gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n483), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n716), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NOR2_X1   g528(.A1(new_n716), .A2(new_n462), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g530(.A1(new_n669), .A2(new_n671), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n541), .A3(new_n579), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n652), .ZN(new_n734));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734), .B2(new_n543), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n541), .A2(new_n579), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n488), .A2(new_n660), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(KEYINPUT108), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n741), .A2(new_n583), .A3(new_n544), .A4(new_n652), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n735), .A2(new_n742), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n734), .B2(new_n285), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n741), .A2(new_n584), .A3(new_n448), .A4(new_n652), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT52), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT109), .B1(new_n734), .B2(new_n285), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n749), .A3(new_n448), .A4(new_n652), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n748), .A2(G92gat), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(new_n751), .B2(new_n753), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n734), .B2(new_n689), .ZN(new_n755));
  INV_X1    g554(.A(G99gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n686), .A2(new_n612), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(G1338gat));
  INV_X1    g558(.A(G106gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n612), .A2(new_n462), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n741), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n736), .B(new_n761), .C1(new_n669), .C2(new_n671), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT53), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n762), .A2(KEYINPUT53), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n760), .B1(new_n763), .B2(KEYINPUT110), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT110), .B2(new_n763), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(G1339gat));
  XOR2_X1   g571(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n773));
  NAND4_X1  g572(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n608), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n601), .A2(KEYINPUT54), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n600), .B1(new_n598), .B2(new_n599), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n609), .B1(new_n779), .B2(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n601), .A2(KEYINPUT54), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n608), .B(new_n774), .C1(new_n781), .C2(new_n777), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(KEYINPUT113), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT113), .B1(new_n782), .B2(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n521), .A2(new_n522), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n525), .A2(new_n526), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n536), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n660), .A2(new_n540), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n782), .A2(new_n783), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n784), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n540), .A2(new_n790), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n630), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n796), .A2(new_n798), .A3(new_n799), .A4(new_n780), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n541), .A3(new_n780), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n612), .A2(new_n797), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n660), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n658), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n631), .A2(new_n541), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n379), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(new_n544), .A3(new_n285), .A4(new_n483), .ZN(new_n810));
  OAI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n710), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n541), .A2(new_n295), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT115), .Z(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n810), .B2(new_n813), .ZN(G1340gat));
  NOR2_X1   g613(.A1(new_n810), .A2(new_n612), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(new_n293), .ZN(G1341gat));
  OAI21_X1  g615(.A(G127gat), .B1(new_n810), .B2(new_n658), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n579), .A2(new_n286), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n810), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT116), .ZN(G1342gat));
  AOI211_X1 g619(.A(new_n630), .B(new_n810), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n821));
  NOR2_X1   g620(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1343gat));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n462), .B1(new_n806), .B2(new_n808), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n780), .A2(new_n793), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n803), .B1(new_n828), .B2(new_n541), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n792), .B(new_n800), .C1(new_n829), .C2(new_n660), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n807), .B1(new_n830), .B2(new_n711), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT57), .B1(new_n831), .B2(new_n462), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n645), .A2(new_n543), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n448), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n827), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(new_n710), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n335), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  INV_X1    g638(.A(new_n825), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n834), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n710), .A2(G141gat), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n840), .B2(new_n834), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n842), .A2(new_n285), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n838), .A2(new_n839), .A3(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n710), .A2(G141gat), .A3(new_n448), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n839), .B1(new_n838), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n824), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n838), .A2(new_n839), .A3(new_n846), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n335), .B1(new_n841), .B2(new_n848), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n852), .B(KEYINPUT118), .C1(new_n839), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(G1344gat));
  NAND3_X1  g654(.A1(new_n842), .A2(new_n285), .A3(new_n845), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n856), .B2(new_n612), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n333), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n836), .A2(KEYINPUT59), .A3(new_n612), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n806), .A2(new_n808), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n379), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n631), .A2(KEYINPUT120), .A3(new_n541), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT120), .B1(new_n631), .B2(new_n541), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n829), .A2(new_n660), .B1(new_n787), .B2(new_n791), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n711), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n826), .B1(new_n867), .B2(new_n462), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n860), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT119), .B1(new_n825), .B2(KEYINPUT57), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n871), .A2(new_n652), .A3(new_n835), .ZN(new_n872));
  NAND2_X1  g671(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n858), .B(new_n859), .C1(new_n872), .C2(new_n873), .ZN(G1345gat));
  OAI21_X1  g673(.A(G155gat), .B1(new_n836), .B2(new_n658), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n579), .A2(new_n337), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n856), .B2(new_n876), .ZN(G1346gat));
  OR2_X1    g676(.A1(new_n836), .A2(new_n630), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n338), .B1(new_n878), .B2(KEYINPUT121), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(KEYINPUT121), .B2(new_n878), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n660), .A2(new_n338), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n856), .B2(new_n881), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n544), .A2(new_n285), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n809), .A2(new_n483), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n710), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT122), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n861), .A2(new_n543), .A3(new_n448), .A4(new_n380), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n541), .A2(new_n218), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G1348gat));
  OAI21_X1  g688(.A(new_n219), .B1(new_n887), .B2(new_n612), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT123), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n809), .A2(G176gat), .A3(new_n757), .A4(new_n883), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(G1349gat));
  INV_X1    g692(.A(new_n224), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n887), .A2(new_n894), .A3(new_n711), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n884), .A2(new_n658), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G183gat), .ZN(new_n897));
  XOR2_X1   g696(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(G1350gat));
  NOR3_X1   g698(.A1(new_n887), .A2(G190gat), .A3(new_n630), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT125), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n225), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n884), .B2(new_n630), .ZN(new_n903));
  NOR2_X1   g702(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(G1351gat));
  NOR3_X1   g706(.A1(new_n645), .A2(new_n544), .A3(new_n285), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n825), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n541), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n871), .A2(new_n908), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n541), .A2(G197gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  OAI21_X1  g714(.A(G204gat), .B1(new_n912), .B2(new_n612), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n909), .A2(G204gat), .A3(new_n612), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1353gat));
  OR3_X1    g718(.A1(new_n909), .A2(G211gat), .A3(new_n711), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n579), .B(new_n908), .C1(new_n869), .C2(new_n870), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT127), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n926), .B(new_n920), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n912), .B2(new_n630), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n630), .A2(G218gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n909), .B2(new_n930), .ZN(G1355gat));
endmodule


