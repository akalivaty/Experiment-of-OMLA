//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n523, new_n524, new_n525, new_n526, new_n527, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n538,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT64), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT65), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n470), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n462), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT66), .Z(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n463), .A2(G138), .A3(new_n462), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n468), .A2(new_n470), .A3(G126), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n462), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT4), .A4(G138), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n498), .A3(new_n500), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n504), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  AOI22_X1  g087(.A1(new_n505), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n498), .A2(new_n500), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n508), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n515), .B1(G51), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT7), .Z(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(G286));
  INV_X1    g096(.A(G286), .ZN(G168));
  AOI22_X1  g097(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n503), .ZN(new_n524));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n506), .A2(new_n525), .B1(new_n508), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n524), .A2(new_n527), .ZN(G301));
  INV_X1    g103(.A(G301), .ZN(G171));
  AOI22_X1  g104(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n503), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT67), .B(G81), .Z(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n506), .A2(new_n532), .B1(new_n508), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(new_n536));
  XOR2_X1   g111(.A(new_n536), .B(KEYINPUT68), .Z(G153));
  AND3_X1   g112(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G36), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G188));
  NAND3_X1  g117(.A1(new_n498), .A2(new_n500), .A3(G65), .ZN(new_n543));
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(KEYINPUT70), .A3(new_n544), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(G651), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n501), .A2(G91), .A3(new_n505), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(KEYINPUT69), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n553), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n505), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n549), .A2(new_n550), .A3(new_n557), .ZN(G299));
  OAI21_X1  g133(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n501), .A2(G87), .A3(new_n505), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G288));
  INV_X1    g138(.A(G86), .ZN(new_n564));
  INV_X1    g139(.A(G48), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n506), .A2(new_n564), .B1(new_n508), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n514), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(KEYINPUT71), .A3(G651), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n567), .A2(new_n573), .A3(new_n574), .ZN(G305));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n506), .A2(new_n576), .B1(new_n508), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT72), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n579), .A2(KEYINPUT72), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n581), .A2(new_n582), .B1(new_n503), .B2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n514), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(G54), .A2(new_n516), .B1(new_n587), .B2(G651), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n506), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT10), .B1(new_n506), .B2(new_n589), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G171), .B2(new_n593), .ZN(G284));
  OAI21_X1  g170(.A(new_n594), .B1(G171), .B2(new_n593), .ZN(G321));
  NAND2_X1  g171(.A1(G299), .A2(new_n593), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G168), .B2(new_n593), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(G168), .B2(new_n593), .ZN(G280));
  INV_X1    g174(.A(new_n592), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  INV_X1    g177(.A(new_n535), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n593), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n592), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n593), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g182(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT73), .B(G2100), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n476), .A2(G123), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n478), .A2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n612), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2435), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2438), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT75), .B(G2443), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n625), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G1341), .B(G1348), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n634), .A2(G14), .ZN(G401));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2072), .B(G2078), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n637), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT77), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(KEYINPUT78), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n644), .B1(new_n647), .B2(new_n641), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n640), .A2(new_n642), .A3(new_n636), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n647), .A2(new_n641), .A3(new_n636), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n618), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n656), .A2(new_n657), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n661), .A3(new_n658), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n667), .C1(new_n661), .C2(new_n666), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(G1986), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT22), .B(G1981), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  INV_X1    g250(.A(G29), .ZN(new_n676));
  NOR2_X1   g251(.A1(G162), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(G35), .ZN(new_n678));
  OAI21_X1  g253(.A(KEYINPUT95), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(KEYINPUT95), .B2(new_n678), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT29), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n676), .A2(G26), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n684));
  INV_X1    g259(.A(G104), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n462), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT89), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n476), .A2(G128), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n478), .A2(G140), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT90), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n683), .B1(new_n691), .B2(G29), .ZN(new_n692));
  MUX2_X1   g267(.A(new_n683), .B(new_n692), .S(KEYINPUT28), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2067), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT87), .B1(G4), .B2(G16), .ZN(new_n695));
  OR3_X1    g270(.A1(KEYINPUT87), .A2(G4), .A3(G16), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n696), .C1(new_n592), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1348), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(G19), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n535), .B2(new_n697), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT88), .B(G1341), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n694), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n676), .A2(G33), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT25), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n478), .A2(G139), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n708), .B(new_n709), .C1(new_n462), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT93), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n706), .B1(new_n713), .B2(new_n676), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2072), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G21), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G168), .B2(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1966), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G28), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(G28), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n721), .A3(new_n676), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n718), .B(new_n722), .C1(new_n676), .C2(new_n617), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G11), .ZN(new_n724));
  NOR2_X1   g299(.A1(G5), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G171), .B2(G16), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n724), .B1(new_n726), .B2(G1961), .C1(new_n717), .C2(G1966), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n478), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n476), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  NAND4_X1  g307(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G32), .B(new_n733), .S(G29), .Z(new_n734));
  XOR2_X1   g309(.A(KEYINPUT27), .B(G1996), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n723), .A2(new_n727), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n676), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n676), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G299), .A2(G16), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n744));
  INV_X1    g319(.A(G20), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G16), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1956), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n737), .A2(new_n741), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n705), .A2(new_n715), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G25), .A2(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n476), .A2(G119), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n478), .A2(G131), .ZN(new_n753));
  NOR2_X1   g328(.A1(G95), .A2(G2105), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT82), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT35), .B(G1991), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n697), .A2(G22), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G166), .B2(new_n697), .ZN(new_n764));
  INV_X1    g339(.A(G1971), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G6), .B(G305), .S(G16), .Z(new_n767));
  XOR2_X1   g342(.A(KEYINPUT32), .B(G1981), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n697), .A2(G23), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n562), .B2(new_n697), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT33), .B(G1976), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT84), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n771), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n766), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G24), .ZN(new_n776));
  XNOR2_X1  g351(.A(G290), .B(KEYINPUT83), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1986), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n762), .B1(KEYINPUT34), .B2(new_n775), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT85), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n775), .A2(KEYINPUT34), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(KEYINPUT86), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n682), .B(new_n750), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(KEYINPUT24), .A2(G34), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT24), .A2(G34), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n791), .A2(new_n676), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G160), .B2(new_n676), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT94), .B(G2084), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n726), .A2(G1961), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n790), .A2(new_n796), .A3(new_n798), .ZN(G311));
  INV_X1    g374(.A(new_n750), .ZN(new_n800));
  INV_X1    g375(.A(new_n789), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n785), .A2(new_n787), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n796), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n803), .A2(new_n804), .A3(new_n797), .A4(new_n682), .ZN(G150));
  AOI22_X1  g380(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n503), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n506), .A2(new_n808), .B1(new_n508), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n592), .A2(new_n601), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT39), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n812), .A2(new_n535), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n603), .A2(new_n811), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n822), .B2(G860), .ZN(G145));
  NAND2_X1  g398(.A1(new_n476), .A2(G130), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n478), .A2(G142), .ZN(new_n825));
  NOR2_X1   g400(.A1(G106), .A2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n756), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n483), .B(G160), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n617), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n495), .B(new_n733), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n691), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n712), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n713), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n834), .A2(new_n842), .A3(new_n840), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n609), .B(KEYINPUT100), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n847), .B1(new_n844), .B2(new_n845), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n830), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(new_n829), .A3(new_n848), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT40), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n851), .A2(new_n853), .A3(new_n857), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(G395));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n860));
  XNOR2_X1  g435(.A(G303), .B(G288), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G290), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G305), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(KEYINPUT42), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n866), .B2(KEYINPUT42), .ZN(new_n867));
  XOR2_X1   g442(.A(G299), .B(new_n592), .Z(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(KEYINPUT41), .B2(new_n869), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n821), .B(new_n605), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n873), .B2(new_n869), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n867), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G868), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n811), .A2(G868), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n860), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI211_X1 g455(.A(KEYINPUT103), .B(new_n878), .C1(new_n876), .C2(G868), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(G295));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n879), .ZN(G331));
  XNOR2_X1  g458(.A(new_n821), .B(G301), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G168), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(new_n872), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n869), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n888), .B2(new_n866), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n866), .B2(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n868), .A2(new_n870), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n885), .B(new_n893), .C1(KEYINPUT41), .C2(new_n868), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  INV_X1    g472(.A(new_n866), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n899), .A2(KEYINPUT43), .A3(new_n889), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT44), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n891), .A3(new_n889), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(KEYINPUT44), .B2(new_n904), .ZN(G397));
  INV_X1    g480(.A(G1384), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n495), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G160), .A2(G40), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n691), .B(G2067), .Z(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n733), .B(G1996), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n912), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n756), .B(new_n761), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR3_X1    g494(.A1(new_n917), .A2(G1986), .A3(G290), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT48), .Z(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n912), .B1(new_n914), .B2(new_n733), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n917), .B2(G1996), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n917), .A2(new_n924), .A3(G1996), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT47), .Z(new_n928));
  NAND3_X1  g503(.A1(new_n916), .A2(new_n761), .A3(new_n758), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(G2067), .B2(new_n691), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n922), .B(new_n928), .C1(new_n912), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G299), .A2(KEYINPUT113), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n549), .A2(new_n933), .A3(new_n550), .A4(new_n557), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n932), .A2(KEYINPUT57), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT57), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT114), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n934), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT57), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(KEYINPUT57), .A3(new_n934), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  AND4_X1   g519(.A1(KEYINPUT112), .A2(new_n495), .A3(new_n944), .A4(new_n906), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n490), .B2(new_n494), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT112), .B1(new_n946), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n949));
  AOI21_X1  g524(.A(new_n911), .B1(new_n907), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G1956), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G40), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n466), .A2(new_n952), .A3(new_n473), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT56), .B(G2072), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n910), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n937), .A2(new_n943), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT115), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n907), .B2(KEYINPUT50), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n946), .A2(KEYINPUT112), .A3(new_n944), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n962), .A2(new_n950), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n956), .B1(new_n964), .B2(G1956), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(KEYINPUT115), .C1(new_n943), .C2(new_n937), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n946), .A2(new_n953), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(G2067), .ZN(new_n969));
  INV_X1    g544(.A(new_n949), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n911), .B1(new_n946), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n907), .A2(KEYINPUT50), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1348), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n967), .B1(new_n592), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n935), .A2(new_n936), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n956), .C1(new_n964), .C2(G1956), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n910), .A2(new_n953), .A3(new_n954), .ZN(new_n980));
  INV_X1    g555(.A(new_n968), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT58), .B(G1341), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n980), .A2(G1996), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n535), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT59), .Z(new_n985));
  OAI21_X1  g560(.A(new_n965), .B1(new_n935), .B2(new_n936), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT61), .B1(new_n986), .B2(new_n978), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT116), .B1(new_n967), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n992), .B(new_n989), .C1(new_n960), .C2(new_n966), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT60), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n969), .C1(new_n973), .C2(new_n974), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT118), .B1(new_n996), .B2(new_n592), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT117), .A3(new_n592), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n975), .A2(KEYINPUT60), .A3(new_n592), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n969), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n971), .A2(new_n972), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT60), .B(new_n1002), .C1(new_n1003), .C2(G1348), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n600), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .A4(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n975), .A2(KEYINPUT60), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT119), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1011), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n979), .B1(new_n994), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  AOI221_X4 g590(.A(new_n1015), .B1(new_n562), .B2(G1976), .C1(new_n946), .C2(new_n953), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n562), .A2(G1976), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1016), .A2(KEYINPUT109), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n562), .A2(G1976), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n968), .A2(new_n1017), .A3(G8), .A4(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n567), .A2(new_n573), .A3(new_n1026), .A4(new_n574), .ZN(new_n1027));
  INV_X1    g602(.A(new_n571), .ZN(new_n1028));
  OAI21_X1  g603(.A(G1981), .B1(new_n1028), .B2(new_n566), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT111), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n981), .A2(new_n1015), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1036), .A3(new_n1031), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n968), .A2(G8), .A3(new_n1022), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT108), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n968), .A2(new_n1041), .A3(G8), .A4(new_n1022), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(KEYINPUT52), .A3(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1025), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT55), .Z(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n962), .A2(new_n950), .A3(new_n1048), .A4(new_n963), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n954), .A2(new_n953), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n946), .A2(new_n908), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n765), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1047), .B1(new_n1053), .B2(new_n1015), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1052), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n973), .A2(G2090), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1046), .B(G8), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1044), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1044), .A2(new_n1054), .A3(KEYINPUT124), .A4(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n980), .B2(G2078), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT122), .ZN(new_n1065));
  INV_X1    g640(.A(new_n485), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n486), .A2(new_n487), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G2105), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(KEYINPUT4), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n906), .B(new_n908), .C1(new_n1069), .C2(new_n493), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n953), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n1072));
  OR4_X1    g647(.A1(new_n1063), .A2(new_n1071), .A3(G2078), .A4(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1003), .A2(G1961), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n1063), .C1(new_n980), .C2(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1065), .A2(new_n1073), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(KEYINPUT54), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1063), .B(G2078), .C1(new_n953), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n910), .A3(new_n954), .A4(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1065), .A2(new_n1074), .A3(new_n1076), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(G171), .B2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1065), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(G301), .A4(new_n1073), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT125), .B1(new_n1077), .B2(G171), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1084), .A2(G171), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT54), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1094));
  INV_X1    g669(.A(G2084), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n971), .A2(new_n972), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(G8), .A3(G286), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(G168), .A3(new_n1096), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1015), .A2(KEYINPUT120), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1099), .A2(KEYINPUT51), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT121), .B(new_n1098), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1085), .A2(new_n1092), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1014), .A2(new_n1062), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1099), .A2(KEYINPUT51), .A3(new_n1100), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1098), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1106), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1105), .A2(new_n1117), .A3(new_n1106), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1116), .A2(new_n1078), .A3(new_n1118), .A4(new_n1062), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT126), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1118), .A2(new_n1078), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1122), .A2(KEYINPUT62), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n981), .A2(new_n1015), .A3(new_n1027), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1015), .B(G286), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1047), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1044), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1054), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1057), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1025), .A2(new_n1043), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1134), .A2(new_n1135), .B1(new_n562), .B2(new_n1016), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1038), .ZN(new_n1137));
  OAI221_X1 g712(.A(new_n1127), .B1(new_n1128), .B2(new_n1132), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1108), .A2(new_n1126), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n912), .A2(G1986), .A3(G290), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n920), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT106), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1140), .A2(KEYINPUT127), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT127), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n931), .B1(new_n1145), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g722(.A(new_n460), .B1(new_n902), .B2(new_n903), .ZN(new_n1149));
  NOR2_X1   g723(.A1(G227), .A2(G401), .ZN(new_n1150));
  NAND4_X1  g724(.A1(new_n855), .A2(new_n1149), .A3(new_n674), .A4(new_n1150), .ZN(G225));
  INV_X1    g725(.A(G225), .ZN(G308));
endmodule


