//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n205), .B(new_n209), .C1(new_n210), .C2(new_n208), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT27), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G183gat), .ZN(new_n216));
  AND4_X1   g015(.A1(KEYINPUT28), .A2(new_n207), .A3(new_n216), .A4(new_n205), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT67), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220));
  AOI211_X1 g019(.A(new_n220), .B(new_n217), .C1(new_n211), .C2(new_n213), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(KEYINPUT26), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(KEYINPUT26), .B2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n219), .A2(new_n221), .A3(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n232), .A2(new_n233), .A3(new_n224), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n205), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(new_n229), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n235), .B(KEYINPUT64), .Z(new_n242));
  OAI211_X1 g041(.A(new_n234), .B(KEYINPUT25), .C1(new_n242), .C2(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n231), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G226gat), .A2(G233gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT72), .Z(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n207), .A2(new_n216), .ZN(new_n251));
  AOI21_X1  g050(.A(G190gat), .B1(new_n251), .B2(KEYINPUT65), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n212), .B1(new_n252), .B2(new_n209), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n220), .B1(new_n253), .B2(new_n217), .ZN(new_n254));
  INV_X1    g053(.A(new_n230), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n214), .A2(KEYINPUT67), .A3(new_n218), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n257), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT73), .B1(new_n257), .B2(new_n244), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT29), .ZN(new_n260));
  INV_X1    g059(.A(new_n247), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n250), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  INV_X1    g063(.A(G211gat), .ZN(new_n265));
  INV_X1    g064(.A(G218gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n268), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n231), .B2(new_n245), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n257), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n261), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n248), .B1(new_n246), .B2(KEYINPUT29), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n268), .B(new_n269), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n204), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT30), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G1gat), .B(G29gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G85gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G57gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G113gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n291), .A2(G120gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n288), .B(new_n289), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT69), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(new_n289), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT68), .B(G113gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(new_n303), .B2(new_n290), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n288), .A4(new_n289), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n298), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G155gat), .B(G162gat), .Z(new_n308));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(G155gat), .B2(G162gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G141gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT76), .B(G141gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G148gat), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n313), .A2(new_n318), .A3(KEYINPUT75), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT75), .B1(new_n313), .B2(new_n318), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n319), .A2(new_n320), .A3(new_n310), .ZN(new_n321));
  INV_X1    g120(.A(new_n308), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(new_n318), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n310), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n318), .A3(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(new_n308), .B1(new_n315), .B2(new_n311), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n331), .A2(new_n302), .A3(new_n298), .A4(new_n306), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT5), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n307), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n316), .B(new_n344), .C1(new_n321), .C2(new_n322), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n307), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n344), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT4), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n335), .B1(new_n348), .B2(new_n332), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n332), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n341), .A2(new_n342), .ZN(new_n355));
  AOI211_X1 g154(.A(new_n352), .B(new_n354), .C1(new_n355), .C2(new_n348), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n287), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n343), .ZN(new_n358));
  INV_X1    g157(.A(new_n337), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n354), .B1(new_n355), .B2(new_n348), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n351), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n286), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(KEYINPUT6), .A3(new_n287), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n272), .A2(new_n279), .A3(new_n204), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n274), .A2(new_n370), .A3(new_n275), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n249), .B1(new_n371), .B2(new_n247), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n279), .B1(new_n372), .B2(new_n278), .ZN(new_n373));
  INV_X1    g172(.A(new_n204), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT74), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n282), .A2(new_n368), .A3(new_n369), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT31), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT78), .B(G50gat), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT79), .B1(new_n278), .B2(KEYINPUT29), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n271), .A2(new_n385), .A3(new_n370), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n344), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n383), .B1(new_n387), .B2(new_n323), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n345), .A2(new_n370), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT80), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n345), .A2(new_n391), .A3(new_n370), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n278), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n278), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n271), .B2(new_n370), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n341), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n383), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n394), .B2(new_n398), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT81), .B(new_n382), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G22gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n382), .A2(KEYINPUT81), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n406), .C1(new_n382), .C2(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n378), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n257), .A2(new_n342), .A3(new_n244), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n342), .B1(new_n257), .B2(new_n244), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n257), .A2(new_n244), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n307), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n411), .B1(new_n422), .B2(new_n413), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n417), .B(new_n420), .C1(KEYINPUT33), .C2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n423), .B2(KEYINPUT33), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT32), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n411), .A3(new_n413), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT34), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n411), .B2(KEYINPUT70), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n422), .A2(new_n411), .A3(new_n413), .A4(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n432), .A2(KEYINPUT71), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT71), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n424), .B(new_n428), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(KEYINPUT71), .A3(new_n434), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n425), .A2(new_n427), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n413), .ZN(new_n440));
  AOI221_X4 g239(.A(new_n426), .B1(KEYINPUT33), .B2(new_n420), .C1(new_n440), .C2(new_n412), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT36), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n282), .A2(new_n369), .A3(new_n377), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT84), .B1(new_n350), .B2(new_n356), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n360), .A2(new_n447), .A3(new_n362), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n286), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n324), .A2(new_n332), .A3(new_n334), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n450), .B2(KEYINPUT82), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n453), .C1(new_n361), .C2(new_n334), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n361), .A2(new_n334), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n286), .B(new_n454), .C1(new_n455), .C2(KEYINPUT39), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT40), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n449), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n409), .B1(new_n445), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT37), .B(new_n279), .C1(new_n372), .C2(new_n278), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n204), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n373), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n465), .B1(new_n464), .B2(new_n204), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT38), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n366), .A2(KEYINPUT6), .A3(new_n287), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n363), .A2(new_n364), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n449), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n276), .A2(new_n277), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n271), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n477), .B(KEYINPUT37), .C1(new_n262), .C2(new_n271), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n468), .A2(new_n478), .A3(new_n479), .A4(new_n204), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n471), .A2(new_n475), .A3(new_n375), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n444), .B1(new_n463), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n474), .A2(new_n282), .A3(new_n369), .A4(new_n377), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n437), .A2(new_n408), .A3(new_n442), .A4(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT86), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n376), .B1(new_n375), .B2(KEYINPUT74), .ZN(new_n487));
  AOI211_X1 g286(.A(new_n281), .B(KEYINPUT30), .C1(new_n373), .C2(new_n374), .ZN(new_n488));
  INV_X1    g287(.A(new_n369), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  AND4_X1   g290(.A1(new_n484), .A2(new_n437), .A3(new_n408), .A4(new_n442), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n474), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n443), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n408), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT35), .B1(new_n496), .B2(new_n378), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n410), .A2(new_n482), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502));
  XNOR2_X1  g301(.A(G57gat), .B(G64gat), .ZN(new_n503));
  INV_X1    g302(.A(G71gat), .ZN(new_n504));
  INV_X1    g303(.A(G78gat), .ZN(new_n505));
  OAI221_X1 g304(.A(new_n501), .B1(new_n502), .B2(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(KEYINPUT91), .A2(G64gat), .ZN(new_n507));
  INV_X1    g306(.A(G57gat), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n508), .A2(G64gat), .ZN(new_n509));
  OAI221_X1 g308(.A(new_n507), .B1(KEYINPUT92), .B2(new_n508), .C1(new_n509), .C2(KEYINPUT91), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT92), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n499), .A2(KEYINPUT9), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n504), .B2(new_n505), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT21), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(new_n265), .ZN(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n517), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n525), .A2(new_n527), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(G1gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT89), .ZN(new_n533));
  AOI21_X1  g332(.A(G8gat), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n532), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n516), .B2(new_n515), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(new_n206), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n536), .B(G183gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G127gat), .B(G155gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT95), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n539), .B2(new_n542), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n523), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G43gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n554), .A2(G50gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(G50gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT15), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT87), .B(G50gat), .Z(new_n559));
  OAI21_X1  g358(.A(new_n555), .B1(new_n559), .B2(G43gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G29gat), .ZN(new_n563));
  INV_X1    g362(.A(G36gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT14), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n565), .B(new_n567), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n557), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT17), .ZN(new_n572));
  OR2_X1    g371(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n573));
  NAND2_X1  g372(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n573), .A2(G85gat), .A3(G92gat), .A4(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(KEYINPUT8), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n575), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n575), .A2(new_n582), .A3(new_n584), .A4(new_n578), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(KEYINPUT97), .A3(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n572), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n571), .A2(new_n591), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n553), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n597), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n552), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n539), .A2(new_n542), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n544), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n522), .A3(new_n546), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n549), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n498), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n572), .A2(new_n535), .ZN(new_n610));
  INV_X1    g409(.A(new_n571), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n611), .A2(new_n535), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n611), .B(new_n535), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n613), .B(KEYINPUT13), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n612), .A4(new_n613), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622));
  INV_X1    g421(.A(G197gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT11), .B(G169gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n616), .A2(new_n627), .A3(new_n619), .A4(new_n620), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n506), .A2(new_n514), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n591), .A2(new_n632), .A3(KEYINPUT10), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n588), .B1(new_n586), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT99), .B1(new_n583), .B2(new_n585), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n515), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n591), .B2(new_n632), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n515), .A2(new_n589), .A3(KEYINPUT98), .A4(new_n590), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n641), .A2(KEYINPUT100), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT100), .B1(new_n641), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n633), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT101), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n648), .B(new_n633), .C1(new_n643), .C2(new_n644), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n641), .A2(new_n647), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT102), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n650), .A2(new_n658), .A3(new_n651), .A4(new_n655), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n631), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n647), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n651), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n654), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n609), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n368), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n526), .ZN(G1324gat));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n490), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n668), .B(KEYINPUT103), .Z(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(G8gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n669), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(new_n665), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n677), .A2(G15gat), .A3(new_n444), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n677), .B2(new_n495), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n408), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  OAI21_X1  g483(.A(KEYINPUT44), .B1(new_n498), .B2(new_n604), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n463), .A2(new_n481), .ZN(new_n686));
  INV_X1    g485(.A(new_n444), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n410), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n378), .A2(KEYINPUT106), .A3(new_n409), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n494), .A2(new_n497), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  INV_X1    g493(.A(new_n604), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n685), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n657), .A2(new_n659), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n549), .A2(new_n607), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n629), .A2(new_n630), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n663), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT105), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT107), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n705), .B(new_n702), .C1(new_n685), .C2(new_n696), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n368), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n498), .A2(new_n604), .A3(new_n701), .ZN(new_n709));
  INV_X1    g508(.A(new_n368), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n563), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(G1328gat));
  OAI21_X1  g512(.A(G36gat), .B1(new_n707), .B2(new_n490), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n709), .A2(new_n564), .A3(new_n445), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT46), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1329gat));
  AOI211_X1 g516(.A(KEYINPUT44), .B(new_n604), .C1(new_n691), .C2(new_n692), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n445), .A2(new_n462), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n408), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n466), .A2(new_n468), .ZN(new_n721));
  INV_X1    g520(.A(new_n470), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n479), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n447), .B1(new_n360), .B2(new_n362), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n350), .A2(KEYINPUT84), .A3(new_n356), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n287), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n473), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(new_n375), .A3(new_n480), .A4(new_n472), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n410), .B(new_n687), .C1(new_n720), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n692), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n694), .B1(new_n732), .B2(new_n695), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n703), .B1(new_n718), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G43gat), .B1(new_n734), .B2(new_n687), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n709), .A2(new_n554), .A3(new_n495), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(KEYINPUT47), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n736), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n444), .B1(new_n704), .B2(new_n706), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n705), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n697), .A2(KEYINPUT107), .A3(new_n703), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n408), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT108), .B1(new_n744), .B2(new_n559), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n709), .A2(new_n559), .A3(new_n409), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n409), .B1(new_n704), .B2(new_n706), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  INV_X1    g547(.A(new_n559), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n745), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n734), .B2(new_n408), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(KEYINPUT48), .A3(new_n746), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1331gat));
  NOR2_X1   g555(.A1(new_n608), .A2(new_n700), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n693), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n698), .A2(new_n663), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n368), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n508), .ZN(G1332gat));
  AOI211_X1 g561(.A(new_n490), .B(new_n760), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n760), .B2(new_n687), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n758), .A2(new_n504), .A3(new_n495), .A4(new_n759), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g568(.A1(new_n760), .A2(new_n408), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(new_n505), .ZN(G1335gat));
  INV_X1    g570(.A(new_n699), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n700), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n693), .A2(new_n695), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT51), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n576), .A4(new_n759), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n773), .A2(new_n759), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT109), .Z(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n685), .B2(new_n696), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n710), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n779), .A2(new_n368), .B1(new_n576), .B2(new_n783), .ZN(G1336gat));
  AND2_X1   g583(.A1(new_n782), .A2(new_n445), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n577), .A3(new_n445), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT111), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n785), .A2(new_n577), .B1(new_n775), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n777), .A2(new_n778), .A3(new_n790), .A4(new_n759), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n782), .A2(new_n444), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n791), .A2(new_n443), .B1(new_n790), .B2(new_n792), .ZN(G1338gat));
  AND2_X1   g592(.A1(new_n782), .A2(new_n409), .ZN(new_n794));
  INV_X1    g593(.A(G106gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n759), .A2(new_n795), .A3(new_n409), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT112), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n795), .B1(new_n775), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g598(.A1(new_n698), .A2(new_n663), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n757), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT113), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n613), .B1(new_n610), .B2(new_n612), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n617), .A2(new_n618), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n626), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n630), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n759), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n645), .A2(new_n813), .A3(new_n647), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n814), .A2(new_n815), .A3(new_n654), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n814), .B2(new_n654), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n645), .A2(new_n647), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n812), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n822), .B(KEYINPUT55), .C1(new_n816), .C2(new_n817), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(new_n698), .A3(new_n700), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n695), .B1(new_n811), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n821), .A2(new_n698), .A3(new_n695), .A4(new_n823), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n809), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n699), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n368), .B1(new_n802), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n496), .A2(new_n445), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n631), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n631), .A2(new_n303), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT116), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n832), .B2(new_n835), .ZN(G1340gat));
  NOR2_X1   g635(.A1(new_n832), .A2(new_n800), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n290), .A2(KEYINPUT117), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n290), .A2(KEYINPUT117), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n837), .B2(new_n839), .ZN(G1341gat));
  NAND2_X1  g640(.A1(new_n831), .A2(new_n772), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g642(.A1(new_n831), .A2(new_n695), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n845));
  XOR2_X1   g644(.A(KEYINPUT56), .B(G134gat), .Z(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(G1343gat));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n811), .A2(new_n824), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n604), .ZN(new_n850));
  INV_X1    g649(.A(new_n827), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n772), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n801), .B(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n848), .B(new_n409), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n444), .A2(new_n368), .A3(new_n445), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n818), .B2(new_n820), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT55), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n857), .B(new_n812), .C1(new_n818), .C2(new_n820), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n660), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n695), .B1(new_n861), .B2(new_n811), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n699), .B1(new_n862), .B2(new_n827), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n408), .B1(new_n863), .B2(new_n802), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n855), .B(new_n856), .C1(new_n864), .C2(new_n848), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n314), .B1(new_n865), .B2(new_n631), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n444), .B1(new_n829), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n710), .B1(new_n852), .B2(new_n854), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n445), .A2(new_n408), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n631), .A2(G141gat), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n869), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n867), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n866), .B(new_n874), .C1(KEYINPUT120), .C2(KEYINPUT58), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(G148gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n759), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n881), .A2(KEYINPUT121), .A3(G148gat), .A4(new_n800), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n408), .B1(new_n802), .B2(new_n828), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(new_n848), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n863), .A2(new_n801), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n848), .A3(new_n409), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n887), .A2(new_n759), .A3(new_n856), .A4(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n885), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n885), .B(G148gat), .C1(new_n865), .C2(new_n800), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n883), .A2(new_n884), .B1(new_n891), .B2(new_n893), .ZN(G1345gat));
  INV_X1    g693(.A(G155gat), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n865), .A2(new_n895), .A3(new_n699), .ZN(new_n896));
  INV_X1    g695(.A(new_n881), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n772), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n895), .ZN(G1346gat));
  INV_X1    g698(.A(G162gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n900), .A3(new_n695), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n865), .A2(new_n604), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(G162gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n901), .B2(new_n905), .ZN(G1347gat));
  AOI21_X1  g705(.A(new_n496), .B1(new_n802), .B2(new_n828), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n490), .A2(new_n710), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n631), .ZN(new_n910));
  XOR2_X1   g709(.A(KEYINPUT123), .B(G169gat), .Z(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1348gat));
  NOR2_X1   g711(.A1(new_n909), .A2(new_n800), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT124), .B(G176gat), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(G1349gat));
  INV_X1    g714(.A(new_n909), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n251), .A3(new_n772), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n206), .B1(new_n909), .B2(new_n699), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n921), .B(new_n922), .Z(G1350gat));
  NAND2_X1  g722(.A1(new_n916), .A2(new_n695), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(G190gat), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n924), .B2(G190gat), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT61), .B(new_n205), .C1(new_n916), .C2(new_n695), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n926), .A2(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1351gat));
  AND2_X1   g730(.A1(new_n887), .A2(new_n889), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n687), .A2(new_n908), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n631), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n886), .A2(new_n934), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n623), .A3(new_n700), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1352gat));
  NAND3_X1  g739(.A1(new_n932), .A2(new_n759), .A3(new_n934), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n937), .A2(G204gat), .A3(new_n800), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT127), .B1(new_n944), .B2(new_n943), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n944), .A2(KEYINPUT127), .A3(new_n943), .ZN(new_n946));
  OAI221_X1 g745(.A(new_n942), .B1(new_n943), .B2(new_n944), .C1(new_n945), .C2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n938), .A2(new_n265), .A3(new_n772), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n887), .A2(new_n772), .A3(new_n889), .A4(new_n934), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n935), .B2(new_n604), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n266), .A3(new_n695), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1355gat));
endmodule


