//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n210), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n202), .A2(new_n203), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  OAI22_X1  g0022(.A1(new_n219), .A2(KEYINPUT0), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT0), .B2(new_n219), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  INV_X1    g0026(.A(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G116), .ZN(new_n228));
  INV_X1    g0028(.A(G270), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n201), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G77), .ZN(new_n232));
  INV_X1    g0032(.A(G244), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n231), .B1(new_n232), .B2(new_n233), .C1(new_n207), .C2(new_n218), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n214), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n225), .A2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  NAND2_X1  g0046(.A1(new_n201), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT67), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT66), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n252), .B(new_n256), .ZN(G351));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n212), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n260), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G13), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n270), .A2(new_n212), .A3(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n258), .A2(new_n259), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n211), .A2(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G50), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n270), .A2(G1), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G20), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(G50), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G223), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n285), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G222), .A3(new_n281), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n287), .B(new_n289), .C1(new_n232), .C2(new_n288), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n259), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n283), .C2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n297), .A2(new_n293), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n295), .B1(new_n298), .B2(G226), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n280), .B1(new_n301), .B2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n309), .A2(new_n261), .B1(new_n212), .B2(new_n232), .ZN(new_n310));
  INV_X1    g0110(.A(new_n267), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n264), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n272), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT70), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n232), .B1(new_n211), .B2(G20), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n273), .A2(new_n315), .B1(new_n232), .B2(new_n271), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n295), .B1(new_n298), .B2(G244), .ZN(new_n319));
  INV_X1    g0119(.A(new_n288), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(G107), .B1(new_n286), .B2(G238), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n288), .A2(G232), .A3(new_n281), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n319), .B1(new_n323), .B2(new_n297), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT71), .B(G200), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n318), .B(new_n327), .C1(new_n328), .C2(new_n324), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n317), .B(new_n331), .C1(G179), .C2(new_n324), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n308), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT9), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n280), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n300), .A2(new_n326), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n292), .A2(G190), .A3(new_n299), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n279), .A2(KEYINPUT9), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT10), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n279), .B(new_n334), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n337), .A4(new_n336), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n288), .A2(G226), .A3(new_n281), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n297), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n349), .B2(new_n348), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n295), .B1(new_n298), .B2(G238), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n351), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g0155(.A(G200), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n353), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT13), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G190), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n263), .A2(G77), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n361), .B1(new_n212), .B2(G68), .C1(new_n201), .C2(new_n311), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n277), .A2(KEYINPUT12), .A3(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT12), .B1(new_n277), .B2(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n203), .B1(new_n211), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n364), .A2(new_n365), .B1(new_n273), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT11), .B1(new_n362), .B2(new_n272), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n356), .A2(new_n360), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(G169), .B1(new_n354), .B2(new_n355), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n358), .A2(new_n359), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(G169), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n358), .A2(G179), .A3(new_n359), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n370), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n368), .A2(KEYINPUT74), .A3(new_n369), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n372), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n273), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n265), .A2(new_n274), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n277), .B2(new_n265), .ZN(new_n389));
  AND2_X1   g0189(.A1(KEYINPUT75), .A2(G33), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT75), .A2(G33), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT3), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(new_n212), .A3(new_n284), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n392), .A2(new_n395), .A3(new_n212), .A4(new_n284), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(G68), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT76), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(G58), .A3(G68), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n401), .A3(new_n221), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n267), .A2(G159), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n397), .A2(new_n406), .A3(KEYINPUT16), .A4(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n409), .A2(new_n272), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  AOI21_X1  g0212(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT7), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT75), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n283), .ZN(new_n417));
  NAND2_X1  g0217(.A1(KEYINPUT75), .A2(G33), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n282), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n284), .A2(new_n413), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n415), .A2(new_n419), .B1(new_n395), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n412), .B1(new_n421), .B2(new_n203), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n395), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT3), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(new_n414), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT78), .A3(G68), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n406), .A2(new_n408), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n411), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n389), .B1(new_n410), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n227), .A2(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G223), .B2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n284), .B2(new_n392), .ZN(new_n433));
  INV_X1    g0233(.A(G87), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n283), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n291), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n295), .B1(new_n298), .B2(G232), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G169), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(G179), .A3(new_n437), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT18), .B1(new_n430), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n389), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n421), .A2(new_n412), .A3(new_n203), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT78), .B1(new_n425), .B2(G68), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n406), .A2(new_n408), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT16), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n409), .A2(new_n272), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  INV_X1    g0251(.A(new_n441), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G200), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n436), .B2(new_n437), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n436), .A2(new_n437), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(G190), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n443), .B(new_n457), .C1(new_n448), .C2(new_n449), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n410), .A2(new_n429), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(KEYINPUT17), .A3(new_n443), .A4(new_n457), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n442), .A2(new_n453), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n344), .A2(new_n386), .A3(new_n464), .ZN(new_n465));
  OR4_X1    g0265(.A1(KEYINPUT22), .A2(new_n320), .A3(G20), .A4(new_n434), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n282), .B1(new_n417), .B2(new_n418), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT3), .A2(G33), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n212), .B(G87), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT22), .B1(new_n469), .B2(KEYINPUT82), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  AOI21_X1  g0271(.A(G20), .B1(new_n392), .B2(new_n284), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(G87), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n466), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n207), .A2(G20), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT23), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n228), .B1(new_n417), .B2(new_n418), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n212), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n475), .B1(new_n474), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n272), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n260), .B(new_n277), .C1(G1), .C2(new_n283), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT25), .B1(new_n271), .B2(new_n207), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n271), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n484), .A2(G107), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n297), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n218), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT75), .B(G33), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G294), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n468), .B1(new_n496), .B2(KEYINPUT3), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n210), .A2(new_n281), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n217), .A2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n495), .B1(new_n502), .B2(new_n291), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT5), .B(G41), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n297), .A3(G274), .A4(new_n490), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT83), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n501), .B1(new_n392), .B2(new_n284), .ZN(new_n507));
  INV_X1    g0307(.A(new_n497), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n291), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n494), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G264), .ZN(new_n511));
  AND4_X1   g0311(.A1(KEYINPUT83), .A2(new_n509), .A3(new_n505), .A4(new_n511), .ZN(new_n512));
  OR3_X1    g0312(.A1(new_n506), .A2(new_n512), .A3(new_n330), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n503), .A2(G179), .A3(new_n505), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n482), .A2(new_n488), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n482), .A2(new_n488), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n328), .B1(new_n506), .B2(new_n512), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n503), .A2(new_n505), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n454), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n515), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n217), .A2(new_n281), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n218), .A2(G1698), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n467), .C2(new_n468), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n320), .A2(G303), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n291), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n505), .B1(new_n494), .B2(new_n229), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n273), .B(G116), .C1(G1), .C2(new_n283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n271), .A2(new_n228), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n258), .A2(new_n259), .B1(G20), .B2(new_n228), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n212), .C1(G33), .C2(new_n206), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT20), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n536), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n532), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n531), .A2(KEYINPUT21), .A3(G169), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n533), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n538), .A2(new_n537), .ZN(new_n543));
  OAI21_X1  g0343(.A(G169), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n297), .B1(new_n525), .B2(new_n526), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n529), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n528), .A2(new_n530), .A3(G190), .ZN(new_n548));
  OAI21_X1  g0348(.A(G200), .B1(new_n545), .B2(new_n529), .ZN(new_n549));
  INV_X1    g0349(.A(new_n539), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(G179), .A3(new_n539), .ZN(new_n552));
  AND4_X1   g0352(.A1(new_n540), .A2(new_n547), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT81), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n233), .A2(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n498), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n555), .A2(new_n233), .ZN(new_n559));
  INV_X1    g0359(.A(new_n285), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n281), .C1(new_n560), .C2(new_n468), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(G1698), .C1(new_n560), .C2(new_n468), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(new_n535), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n297), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n505), .B1(new_n494), .B2(new_n217), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n554), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n392), .A2(new_n284), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT4), .B1(new_n567), .B2(new_n556), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n535), .A3(new_n562), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n291), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n565), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(KEYINPUT81), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n566), .A2(new_n572), .A3(G190), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT79), .B1(new_n271), .B2(new_n206), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n271), .A2(new_n206), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n574), .B(new_n577), .C1(new_n484), .C2(G97), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n421), .A2(new_n207), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT6), .B1(new_n208), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n583), .A2(new_n212), .B1(new_n232), .B2(new_n311), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n272), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n570), .A2(new_n571), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(G200), .ZN(new_n589));
  INV_X1    g0389(.A(new_n535), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n286), .B2(G250), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n557), .B1(new_n392), .B2(new_n284), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n561), .C1(new_n592), .C2(KEYINPUT4), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n565), .B1(new_n593), .B2(new_n291), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n454), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n573), .B(new_n586), .C1(new_n589), .C2(new_n595), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n554), .B(new_n565), .C1(new_n593), .C2(new_n291), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT81), .B1(new_n570), .B2(new_n571), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n330), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n585), .A2(new_n578), .B1(new_n594), .B2(new_n306), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G238), .A2(G1698), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n233), .B2(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n567), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n478), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n297), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n297), .B(G250), .C1(G1), .C2(new_n489), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n490), .A2(G274), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n326), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n309), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n277), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n567), .A2(new_n212), .A3(G68), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n212), .B1(new_n347), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n434), .A2(new_n206), .A3(new_n207), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n261), .B2(new_n206), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n612), .B1(new_n620), .B2(new_n272), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n484), .A2(G87), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n607), .A2(new_n608), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n478), .B1(new_n567), .B2(new_n603), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(G190), .C1(new_n624), .C2(new_n297), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n610), .A2(new_n621), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n330), .B1(new_n606), .B2(new_n609), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n484), .A2(new_n611), .ZN(new_n628));
  INV_X1    g0428(.A(new_n612), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n617), .A2(new_n618), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(G68), .B2(new_n472), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n628), .B(new_n629), .C1(new_n631), .C2(new_n260), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n623), .B(new_n306), .C1(new_n624), .C2(new_n297), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n553), .A2(new_n596), .A3(new_n601), .A4(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n465), .A2(new_n522), .A3(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n308), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n430), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n451), .B1(new_n450), .B2(new_n452), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n332), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n381), .A2(new_n385), .B1(new_n371), .B2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n460), .A2(new_n462), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n641), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n340), .A2(KEYINPUT85), .A3(new_n343), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT85), .B1(new_n340), .B2(new_n343), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n638), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n465), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n596), .A2(new_n601), .A3(new_n635), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n482), .A2(new_n521), .A3(new_n488), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n547), .A2(new_n540), .A3(new_n552), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n652), .B(new_n653), .C1(new_n655), .C2(new_n515), .ZN(new_n656));
  INV_X1    g0456(.A(new_n634), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n599), .A2(new_n600), .A3(new_n634), .A4(new_n626), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n635), .A2(KEYINPUT26), .A3(new_n599), .A4(new_n600), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n650), .B1(new_n651), .B2(new_n664), .ZN(G369));
  NAND2_X1  g0465(.A1(new_n276), .A2(new_n212), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  INV_X1    g0468(.A(G213), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n666), .B2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n550), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT87), .ZN(new_n675));
  MUX2_X1   g0475(.A(new_n655), .B(new_n553), .S(new_n675), .Z(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n522), .B1(new_n517), .B2(new_n673), .ZN(new_n678));
  INV_X1    g0478(.A(new_n515), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n515), .A2(new_n673), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n654), .A2(new_n673), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n522), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(G399));
  NOR2_X1   g0485(.A1(new_n216), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n616), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n222), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n653), .A2(new_n601), .A3(new_n596), .A4(new_n635), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n513), .A2(new_n514), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n654), .B1(new_n516), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n662), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n673), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT88), .B1(new_n695), .B2(new_n673), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT29), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n673), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n656), .B2(new_n662), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n636), .A2(new_n679), .A3(new_n653), .A4(new_n673), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n546), .A2(G179), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n623), .B1(new_n624), .B2(new_n297), .ZN(new_n706));
  AND4_X1   g0506(.A1(new_n519), .A2(new_n705), .A3(new_n588), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n509), .A2(new_n511), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n531), .A2(new_n306), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n566), .A4(new_n572), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n712), .B2(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n699), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n704), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT31), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n714), .B2(new_n699), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n703), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n702), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n270), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n211), .B1(new_n725), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n686), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n677), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n676), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n676), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n259), .B1(G20), .B2(new_n330), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n212), .A2(new_n328), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n306), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n212), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n741), .A2(G322), .B1(new_n745), .B2(G329), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n739), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n746), .B(new_n320), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n212), .B1(new_n743), .B2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(G294), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n212), .A2(new_n306), .A3(new_n454), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n328), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(G190), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G326), .A2(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  INV_X1    g0559(.A(new_n742), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n325), .A2(new_n760), .A3(G179), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n752), .B(new_n758), .C1(new_n759), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n326), .A2(new_n306), .A3(new_n738), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n763), .B1(G303), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n750), .B(KEYINPUT94), .Z(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G97), .ZN(new_n768));
  INV_X1    g0568(.A(new_n755), .ZN(new_n769));
  INV_X1    g0569(.A(new_n756), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n768), .B1(new_n769), .B2(new_n201), .C1(new_n203), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n762), .A2(new_n207), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n288), .B1(new_n748), .B2(new_n232), .C1(new_n202), .C2(new_n740), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n744), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n434), .B2(new_n764), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n737), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n728), .B(KEYINPUT90), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n216), .A2(new_n567), .ZN(new_n781));
  INV_X1    g0581(.A(new_n222), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n489), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n781), .B(new_n783), .C1(new_n251), .C2(new_n489), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n216), .A2(new_n320), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G355), .B1(new_n228), .B2(new_n216), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT91), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n734), .A2(new_n737), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n787), .B2(KEYINPUT91), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n780), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT92), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n779), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n731), .B1(new_n736), .B2(new_n795), .ZN(G396));
  NOR2_X1   g0596(.A1(new_n332), .A2(new_n699), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n699), .A2(new_n317), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n329), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(new_n799), .B2(new_n332), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n733), .ZN(new_n801));
  INV_X1    g0601(.A(new_n737), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n733), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n780), .B1(G77), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G283), .A2(new_n756), .B1(new_n755), .B2(G303), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n762), .A2(new_n434), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n320), .B1(new_n748), .B2(new_n228), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n740), .A2(new_n808), .B1(new_n744), .B2(new_n747), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n765), .A2(G107), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n768), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n748), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G143), .A2(new_n741), .B1(new_n813), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n769), .B2(new_n815), .C1(new_n816), .C2(new_n770), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n498), .B1(G132), .B2(new_n745), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n202), .B2(new_n750), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G68), .B2(new_n761), .ZN(new_n822));
  INV_X1    g0622(.A(new_n765), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n819), .B(new_n822), .C1(new_n201), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n817), .A2(new_n818), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n812), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT96), .Z(new_n827));
  AOI211_X1 g0627(.A(new_n801), .B(new_n804), .C1(new_n827), .C2(new_n737), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n700), .A2(new_n800), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT97), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n800), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n700), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n721), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n728), .B1(new_n721), .B2(new_n832), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  NOR2_X1   g0637(.A1(new_n725), .A2(new_n211), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n717), .A2(new_n719), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n394), .A2(G68), .A3(new_n396), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n411), .B1(new_n428), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(new_n272), .A3(new_n409), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n671), .B1(new_n842), .B2(new_n443), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n463), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n450), .A2(new_n452), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n450), .A2(new_n672), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n458), .ZN(new_n848));
  INV_X1    g0648(.A(new_n458), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n842), .A2(new_n443), .B1(new_n441), .B2(new_n671), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n845), .A2(new_n846), .A3(new_n458), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  INV_X1    g0655(.A(new_n846), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n855), .A2(new_n848), .B1(new_n463), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n853), .B1(new_n857), .B2(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(new_n800), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n380), .B1(new_n373), .B2(new_n376), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n375), .B1(new_n378), .B2(G169), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n385), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n385), .A2(new_n699), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n371), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n385), .B(new_n699), .C1(new_n381), .C2(new_n372), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n859), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n839), .A2(new_n858), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT31), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n704), .B2(new_n715), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n718), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n865), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n800), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n843), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n641), .B2(new_n644), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n848), .A2(new_n851), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT40), .B1(new_n878), .B2(new_n853), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n867), .A2(KEYINPUT40), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n651), .B2(new_n870), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n866), .B1(new_n869), .B2(new_n718), .ZN(new_n882));
  INV_X1    g0682(.A(new_n858), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT40), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n879), .A2(new_n839), .A3(new_n866), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n465), .A3(new_n839), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(new_n887), .A3(G330), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT100), .Z(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n381), .A2(new_n385), .A3(new_n673), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n844), .B2(new_n852), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT39), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT99), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n853), .B(new_n897), .C1(new_n857), .C2(KEYINPUT38), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n895), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n641), .A2(new_n672), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n797), .B1(new_n700), .B2(new_n800), .ZN(new_n903));
  INV_X1    g0703(.A(new_n871), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n878), .A2(new_n853), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n698), .A2(new_n465), .A3(new_n701), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n650), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n838), .B1(new_n890), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n890), .B2(new_n911), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT35), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n228), .B(new_n220), .C1(new_n583), .C2(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n915), .A2(KEYINPUT98), .B1(new_n914), .B2(new_n583), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(KEYINPUT98), .B2(new_n915), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT36), .Z(new_n918));
  NAND4_X1  g0718(.A1(new_n782), .A2(G77), .A3(new_n401), .A4(new_n399), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n247), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n270), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n913), .A2(new_n918), .A3(new_n921), .ZN(G367));
  AOI22_X1  g0722(.A1(new_n756), .A2(G159), .B1(G68), .B2(new_n767), .ZN(new_n923));
  INV_X1    g0723(.A(new_n764), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G58), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n288), .B1(new_n740), .B2(new_n816), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n748), .A2(new_n201), .B1(new_n744), .B2(new_n815), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(G77), .C2(new_n761), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n755), .A2(G143), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n923), .A2(new_n925), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n755), .A2(G311), .B1(G303), .B2(new_n741), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT108), .Z(new_n932));
  NOR2_X1   g0732(.A1(new_n750), .A2(new_n207), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n745), .A2(G317), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n498), .C1(new_n759), .C2(new_n748), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G97), .C2(new_n761), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n932), .B(new_n936), .C1(new_n808), .C2(new_n770), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n228), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n765), .A2(G116), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(KEYINPUT46), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n930), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT109), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT47), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n737), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n673), .B1(new_n621), .B2(new_n622), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n635), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n634), .B2(new_n945), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT101), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n734), .ZN(new_n949));
  INV_X1    g0749(.A(new_n780), .ZN(new_n950));
  INV_X1    g0750(.A(new_n781), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n245), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n789), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n216), .B2(new_n611), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n944), .A2(new_n949), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n684), .A2(new_n682), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n596), .B(new_n601), .C1(new_n586), .C2(new_n673), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n599), .A2(new_n699), .A3(new_n600), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT44), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n684), .A2(new_n682), .A3(new_n961), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n681), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n957), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n964), .A2(new_n967), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT106), .A3(new_n681), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT104), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n681), .B(KEYINPUT105), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n972), .A2(KEYINPUT104), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n684), .B1(new_n680), .B2(new_n683), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n677), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n723), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n974), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n723), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT107), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n686), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n982), .B1(new_n971), .B2(new_n973), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n722), .B1(new_n990), .B2(new_n979), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT107), .B1(new_n991), .B2(new_n987), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n727), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n522), .A2(new_n683), .A3(new_n961), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n601), .B1(new_n679), .B2(new_n959), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n673), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT102), .Z(new_n1000));
  INV_X1    g0800(.A(new_n948), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n970), .A3(new_n961), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT103), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n681), .B2(new_n962), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n956), .B1(new_n993), .B2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n680), .A2(new_n735), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n688), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n785), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(G107), .B2(new_n215), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n241), .A2(new_n489), .ZN(new_n1018));
  AOI211_X1 g0818(.A(G45), .B(new_n1015), .C1(G68), .C2(G77), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n264), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n951), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1017), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n780), .B1(new_n1023), .B2(new_n953), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT110), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G317), .A2(new_n741), .B1(new_n813), .B2(G303), .ZN(new_n1026));
  INV_X1    g0826(.A(G322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n769), .B2(new_n1027), .C1(new_n747), .C2(new_n770), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n924), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n762), .A2(new_n228), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n567), .B(new_n1037), .C1(G326), .C2(new_n745), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G159), .A2(new_n755), .B1(new_n756), .B2(new_n265), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n748), .A2(new_n203), .B1(new_n744), .B2(new_n816), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n498), .B(new_n1041), .C1(G50), .C2(new_n741), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n924), .A2(G77), .B1(G97), .B2(new_n761), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n767), .A2(new_n611), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1025), .B1(new_n1046), .B2(new_n737), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n981), .A2(new_n727), .B1(new_n1014), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n982), .A2(new_n686), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n723), .A2(new_n981), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(G393));
  AOI22_X1  g0851(.A1(new_n971), .A2(new_n973), .B1(new_n970), .B2(new_n969), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n984), .B(new_n686), .C1(new_n983), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n962), .A2(new_n734), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n256), .A2(new_n951), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n789), .B1(new_n206), .B2(new_n215), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n780), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n769), .A2(new_n816), .B1(new_n774), .B2(new_n740), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G143), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n567), .B1(new_n1061), .B2(new_n744), .C1(new_n264), .C2(new_n748), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1062), .B(new_n806), .C1(G68), .C2(new_n924), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n767), .A2(G77), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n756), .A2(G50), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n755), .A2(G317), .B1(G311), .B2(new_n741), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT52), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n772), .B1(G283), .B2(new_n924), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n756), .A2(G303), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n320), .B1(new_n744), .B2(new_n1027), .C1(new_n808), .C2(new_n748), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G116), .B2(new_n751), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1066), .A2(new_n1067), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1057), .B1(new_n1075), .B2(new_n737), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1052), .A2(new_n727), .B1(new_n1054), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1053), .A2(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(new_n898), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n897), .B1(new_n878), .B2(new_n853), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT99), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n891), .B1(new_n903), .B2(new_n904), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n839), .A2(G330), .A3(new_n866), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n883), .A2(new_n892), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n695), .A2(new_n673), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT88), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n673), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n797), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n799), .A2(new_n332), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1086), .B1(new_n1094), .B2(new_n904), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1084), .A2(new_n1085), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1085), .B1(new_n1084), .B2(new_n1095), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n831), .C1(new_n869), .C2(new_n718), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n904), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1094), .A2(new_n1100), .A3(new_n1085), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n800), .C1(new_n869), .C2(new_n718), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n720), .A2(new_n866), .B1(new_n1102), .B2(new_n904), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n903), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n720), .A2(new_n465), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n909), .A2(new_n650), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT112), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n909), .A2(new_n1105), .A3(KEYINPUT112), .A4(new_n650), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n686), .B1(new_n1098), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT113), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1098), .A2(new_n1112), .A3(new_n1110), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1085), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1084), .A2(new_n1095), .A3(new_n1085), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1111), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n741), .A2(G132), .B1(new_n745), .B2(G125), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n761), .A2(G50), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n320), .B1(new_n813), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n767), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n770), .A2(new_n815), .B1(new_n774), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(G128), .C2(new_n755), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n764), .A2(new_n816), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n756), .A2(G107), .B1(G97), .B2(new_n813), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT115), .Z(new_n1135));
  OAI221_X1 g0935(.A(new_n320), .B1(new_n744), .B2(new_n808), .C1(new_n228), .C2(new_n740), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G68), .B2(new_n761), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1064), .B(new_n1137), .C1(new_n769), .C2(new_n759), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G87), .B2(new_n765), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1130), .A2(new_n1133), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n780), .B1(new_n265), .B2(new_n803), .C1(new_n1140), .C2(new_n802), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n899), .A2(new_n900), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n732), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1098), .B2(new_n727), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1121), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  OAI21_X1  g0947(.A(new_n308), .B1(new_n647), .B2(new_n648), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n279), .A2(new_n671), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n308), .B1(new_n279), .B2(new_n671), .C1(new_n647), .C2(new_n648), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n732), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n728), .B1(G50), .B2(new_n803), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n567), .A2(G41), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n283), .A2(new_n296), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT116), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1158), .A2(G50), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT117), .Z(new_n1162));
  OAI22_X1  g0962(.A1(new_n740), .A2(new_n207), .B1(new_n744), .B2(new_n759), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n611), .B2(new_n813), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n924), .A2(G77), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n761), .A2(G58), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1158), .A4(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n770), .A2(new_n206), .B1(new_n203), .B2(new_n1128), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(G116), .C2(new_n755), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1162), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1128), .A2(new_n816), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n756), .A2(G132), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G128), .A2(new_n741), .B1(new_n813), .B2(G137), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n764), .C2(new_n1124), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1173), .B(new_n1176), .C1(G125), .C2(new_n755), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n761), .A2(G159), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n745), .A2(G124), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1160), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1157), .B1(new_n1185), .B2(new_n737), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1156), .A2(KEYINPUT120), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT120), .B1(new_n1156), .B2(new_n1186), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1155), .B1(new_n880), .B2(new_n703), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1155), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n886), .A2(new_n1193), .A3(G330), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1192), .A2(new_n901), .A3(new_n907), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n886), .B2(G330), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n703), .B(new_n1155), .C1(new_n884), .C2(new_n885), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n908), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1198), .A3(KEYINPUT121), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(KEYINPUT121), .B2(new_n1198), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1191), .B1(new_n1200), .B2(new_n726), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1200), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1112), .B1(new_n1098), .B2(new_n1110), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1119), .A2(new_n1096), .A3(new_n1097), .A4(KEYINPUT113), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1204), .B1(new_n1120), .B2(new_n1113), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n686), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1202), .B1(new_n1209), .B2(new_n1214), .ZN(G375));
  INV_X1    g1015(.A(new_n1102), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1085), .B1(new_n1216), .B2(new_n871), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n903), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n726), .B1(new_n1219), .B2(new_n1101), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n780), .B1(G68), .B2(new_n803), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n871), .A2(new_n733), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n288), .B1(new_n745), .B2(G303), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n207), .B2(new_n748), .C1(new_n759), .C2(new_n740), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G77), .B2(new_n761), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G116), .A2(new_n756), .B1(new_n755), .B2(G294), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n765), .A2(G97), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1044), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1166), .A2(new_n567), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT122), .Z(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n774), .B2(new_n823), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G132), .A2(new_n755), .B1(new_n756), .B2(new_n1125), .ZN(new_n1232));
  INV_X1    g1032(.A(G128), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n740), .A2(new_n815), .B1(new_n744), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G150), .B2(new_n813), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1232), .B(new_n1235), .C1(new_n201), .C2(new_n1128), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1221), .B(new_n1222), .C1(new_n737), .C2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT123), .B1(new_n1220), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1104), .B2(new_n727), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT123), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1119), .A2(new_n988), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(G381));
  INV_X1    g1046(.A(new_n956), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n986), .B1(new_n985), .B2(new_n988), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n991), .A2(KEYINPUT107), .A3(new_n987), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n726), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1247), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT124), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n687), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1211), .B1(new_n1210), .B2(new_n1200), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1201), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1146), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1256), .A2(new_n1260), .ZN(G407));
  NOR2_X1   g1061(.A1(new_n669), .A2(G343), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1146), .A3(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G213), .B(new_n1263), .C1(new_n1256), .C2(new_n1260), .ZN(G409));
  XNOR2_X1  g1064(.A(G393), .B(G396), .ZN(new_n1265));
  XOR2_X1   g1065(.A(G390), .B(new_n1265), .Z(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(G387), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G390), .B(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1252), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1196), .A2(new_n908), .A3(new_n1197), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1192), .A2(new_n1194), .B1(new_n901), .B2(new_n907), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n727), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1191), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1121), .A2(new_n1145), .A3(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1203), .A2(new_n1208), .A3(new_n988), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1262), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1244), .B1(KEYINPUT60), .B2(new_n1119), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1204), .A2(KEYINPUT60), .A3(new_n1219), .A4(new_n1101), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n686), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1243), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n836), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1243), .B(G384), .C1(new_n1278), .C2(new_n1280), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1277), .B(new_n1284), .C1(new_n1259), .C2(new_n1146), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G375), .A2(G378), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1288), .A2(KEYINPUT62), .A3(new_n1284), .A4(new_n1277), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1287), .A2(KEYINPUT127), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(new_n1291), .A3(new_n1286), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1262), .ZN(new_n1293));
  INV_X1    g1093(.A(G2897), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1282), .A2(new_n1297), .A3(new_n1283), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1296), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1295), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1259), .A2(new_n1146), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1111), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1305), .A2(new_n1144), .A3(new_n1191), .A4(new_n1273), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1210), .A2(new_n1200), .A3(new_n987), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1293), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1301), .B(new_n1302), .C1(new_n1303), .C2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1292), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1270), .B1(new_n1290), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1308), .B1(G378), .B2(G375), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1313), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1284), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1315), .B1(new_n1285), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1270), .B1(new_n1316), .B2(new_n1285), .ZN(new_n1319));
  AND2_X1   g1119(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1312), .A2(new_n1321), .ZN(G405));
  NAND2_X1  g1122(.A1(new_n1288), .A2(new_n1260), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1323), .A2(new_n1284), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1270), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1284), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


