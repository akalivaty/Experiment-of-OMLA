//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1189, new_n1190, new_n1191;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n463), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n462), .A3(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G101), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n464), .A2(new_n466), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n463), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G102), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n489), .A2(new_n491), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n507), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n504), .A2(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n502), .A2(new_n514), .ZN(G166));
  INV_X1    g090(.A(new_n512), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n507), .A2(new_n509), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n526));
  INV_X1    g101(.A(new_n504), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n526), .B1(new_n525), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n517), .B(new_n519), .C1(new_n529), .C2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n522), .B2(new_n523), .ZN(new_n534));
  AND2_X1   g109(.A1(G77), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n504), .A2(new_n537), .B1(new_n512), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n522), .B2(new_n523), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT70), .B(G81), .Z(new_n548));
  OAI22_X1  g123(.A1(new_n504), .A2(new_n547), .B1(new_n512), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n520), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g138(.A(KEYINPUT71), .B(new_n559), .C1(new_n520), .C2(new_n560), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(new_n564), .A3(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n516), .A2(G91), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n504), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n503), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(G299));
  OR2_X1    g147(.A1(new_n502), .A2(new_n514), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(G49), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n504), .A2(new_n575), .B1(new_n512), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G288));
  OAI211_X1 g154(.A(G48), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n512), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n501), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n501), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n504), .A2(new_n590), .B1(new_n512), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n512), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n527), .A2(G54), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n501), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n595), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n595), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G299), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G168), .B2(new_n606), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(G168), .B2(new_n606), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n603), .B1(new_n610), .B2(G860), .ZN(G148));
  NOR2_X1   g186(.A1(new_n602), .A2(G559), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n612), .A2(KEYINPUT72), .A3(new_n606), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT72), .B1(new_n612), .B2(new_n606), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G868), .C2(new_n552), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g191(.A1(new_n470), .A2(new_n472), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n495), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n478), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n480), .A2(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2443), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT74), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT75), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n639), .A2(new_n642), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(KEYINPUT75), .A3(new_n642), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n645), .A2(new_n646), .A3(G14), .A4(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT17), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(new_n657), .C2(new_n653), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  AOI22_X1  g246(.A1(new_n669), .A2(KEYINPUT20), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n665), .A3(new_n668), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n674), .C1(KEYINPUT20), .C2(new_n669), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT76), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1971), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n683), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT79), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n683), .A2(G6), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n586), .B2(new_n683), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n692), .B(new_n696), .C1(new_n691), .C2(new_n690), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT77), .B(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n478), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n480), .A2(G131), .ZN(new_n702));
  NOR2_X1   g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT78), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n683), .A2(G24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n593), .B2(new_n683), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n697), .B2(KEYINPUT34), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n698), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT80), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT36), .ZN(new_n717));
  INV_X1    g292(.A(new_n699), .ZN(new_n718));
  AOI21_X1  g293(.A(KEYINPUT28), .B1(new_n718), .B2(G26), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n718), .A2(KEYINPUT28), .A3(G26), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n478), .A2(G128), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT81), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G140), .B2(new_n480), .ZN(new_n723));
  OR2_X1    g298(.A1(G104), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n719), .B(new_n720), .C1(new_n726), .C2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2067), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n552), .A2(new_n683), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n683), .B2(G19), .ZN(new_n730));
  INV_X1    g305(.A(G1341), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n718), .A2(G35), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G162), .B2(new_n718), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT29), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n728), .B(new_n732), .C1(G2090), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G2090), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT87), .Z(new_n738));
  NAND2_X1  g313(.A1(G299), .A2(G16), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT88), .B(KEYINPUT23), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n683), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n603), .A2(new_n683), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G4), .B2(new_n683), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n745), .B1(new_n730), .B2(new_n731), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n736), .A2(new_n738), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n683), .A2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G168), .B2(new_n683), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT84), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1966), .ZN(new_n754));
  NAND2_X1  g329(.A1(G171), .A2(G16), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G5), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  NAND2_X1  g334(.A1(G160), .A2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G34), .Z(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n699), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT82), .B1(G29), .B2(G32), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n478), .A2(G129), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n480), .A2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n617), .A2(G105), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  NAND4_X1  g343(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  MUX2_X1   g346(.A(KEYINPUT82), .B(new_n763), .S(new_n771), .Z(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n758), .B1(new_n759), .B2(new_n762), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n490), .A2(G103), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n480), .A2(G139), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n776), .B(new_n777), .C1(new_n462), .C2(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G33), .B(new_n779), .S(G29), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2072), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT30), .B(G28), .Z(new_n782));
  OAI22_X1  g357(.A1(new_n626), .A2(new_n718), .B1(G29), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n762), .B2(new_n759), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n497), .A2(new_n718), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n699), .A2(G27), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n784), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n774), .A2(new_n781), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n756), .A2(new_n757), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT85), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n772), .A2(new_n773), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT83), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n754), .A2(new_n792), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n750), .B1(new_n797), .B2(KEYINPUT86), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(KEYINPUT86), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n717), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n747), .A2(new_n748), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n716), .A2(KEYINPUT36), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(G311));
  INV_X1    g379(.A(new_n803), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n805), .A2(new_n801), .A3(new_n717), .A4(new_n799), .ZN(G150));
  NAND2_X1  g381(.A1(new_n524), .A2(G67), .ZN(new_n807));
  NAND2_X1  g382(.A1(G80), .A2(G543), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n501), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT89), .B(G55), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n504), .A2(new_n810), .B1(new_n512), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(G860), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT90), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT37), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n809), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(new_n551), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n546), .B(new_n550), .C1(new_n809), .C2(new_n812), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT39), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n603), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n815), .B1(new_n823), .B2(G860), .ZN(G145));
  NAND2_X1  g399(.A1(new_n478), .A2(G130), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n480), .A2(G142), .ZN(new_n826));
  NOR2_X1   g401(.A1(G106), .A2(G2105), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n619), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n705), .ZN(new_n831));
  INV_X1    g406(.A(new_n726), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n769), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n769), .B1(new_n723), .B2(new_n725), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n779), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n833), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n837), .B(KEYINPUT91), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n726), .A2(new_n770), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n834), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n843), .A3(G164), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(G164), .B1(new_n840), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n831), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n840), .A2(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n497), .ZN(new_n849));
  INV_X1    g424(.A(new_n831), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(new_n850), .A3(new_n844), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n626), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n847), .A2(new_n851), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n851), .A2(new_n855), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT93), .B(G37), .Z(new_n858));
  OAI221_X1 g433(.A(new_n831), .B1(KEYINPUT94), .B2(new_n854), .C1(new_n845), .C2(new_n846), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g436(.A(new_n586), .B(KEYINPUT97), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n593), .B(G166), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G288), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n864), .A2(G288), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n864), .A2(G288), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n862), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT42), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT98), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n871), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n819), .B(new_n612), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n602), .A2(KEYINPUT95), .A3(G299), .ZN(new_n879));
  OR2_X1    g454(.A1(G299), .A2(KEYINPUT95), .ZN(new_n880));
  NAND2_X1  g455(.A1(G299), .A2(KEYINPUT95), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n603), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n883), .A2(KEYINPUT96), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(KEYINPUT96), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n882), .B2(new_n879), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n878), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n873), .A2(new_n877), .A3(new_n889), .ZN(new_n890));
  OR3_X1    g465(.A1(new_n872), .A2(new_n889), .A3(KEYINPUT98), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(G868), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(G868), .B2(new_n816), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT99), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G295));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n896), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n900));
  NAND3_X1  g475(.A1(G286), .A2(new_n900), .A3(G301), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(G301), .A2(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT100), .B1(new_n536), .B2(new_n540), .ZN(new_n904));
  NOR3_X1   g479(.A1(G286), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n817), .A2(new_n818), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n817), .B2(new_n818), .ZN(new_n908));
  OAI22_X1  g483(.A1(new_n902), .A2(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n903), .ZN(new_n910));
  INV_X1    g485(.A(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(G168), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n819), .A2(KEYINPUT101), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n817), .A2(new_n818), .A3(new_n906), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(new_n901), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n882), .A2(new_n879), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n886), .A2(new_n887), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n871), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  INV_X1    g501(.A(new_n871), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(new_n918), .C1(new_n921), .C2(new_n922), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n899), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n918), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n916), .A2(new_n920), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n871), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n934), .A2(new_n858), .A3(new_n928), .ZN(new_n935));
  OAI221_X1 g510(.A(new_n931), .B1(new_n930), .B2(new_n929), .C1(new_n925), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n934), .A2(new_n928), .A3(new_n925), .A4(new_n858), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n899), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(G397));
  XNOR2_X1  g517(.A(KEYINPUT104), .B(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n497), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(G160), .A2(G40), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G2067), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n726), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n951), .B2(new_n770), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT46), .Z(new_n955));
  NOR2_X1   g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n956), .B(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n769), .B(new_n953), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n709), .A3(new_n706), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n832), .A2(new_n950), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n949), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT125), .Z(new_n964));
  XOR2_X1   g539(.A(new_n708), .B(KEYINPUT105), .Z(new_n965));
  XNOR2_X1  g540(.A(new_n705), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n948), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT48), .Z(new_n970));
  AOI211_X1 g545(.A(new_n958), .B(new_n964), .C1(new_n968), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n582), .A2(KEYINPUT106), .ZN(new_n973));
  INV_X1    g548(.A(new_n585), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n580), .C1(new_n512), .C2(new_n581), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G1981), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n582), .A2(new_n585), .A3(G1981), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n977), .B2(G1981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n980), .B(KEYINPUT49), .C1(new_n979), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n977), .A2(G1981), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT107), .B1(new_n986), .B2(new_n981), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(KEYINPUT108), .A3(KEYINPUT49), .A4(new_n980), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  INV_X1    g564(.A(new_n980), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n982), .A2(new_n979), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  INV_X1    g568(.A(new_n487), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n495), .B2(G126), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n491), .B1(new_n995), .B2(new_n462), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n494), .A2(new_n496), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(new_n947), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n985), .A2(new_n988), .A3(new_n992), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1003), .B2(G288), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n688), .A2(G1976), .ZN(new_n1005));
  OR3_X1    g580(.A1(new_n1004), .A2(KEYINPUT52), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1002), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G303), .A2(G8), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n469), .A2(new_n475), .A3(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT45), .B(new_n943), .C1(new_n996), .C2(new_n997), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n494), .A2(new_n496), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n488), .A2(G2105), .B1(G102), .B2(new_n490), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1014), .C1(new_n1017), .C2(KEYINPUT45), .ZN(new_n1018));
  INV_X1    g593(.A(G1971), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(G2090), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n497), .A2(new_n1023), .A3(new_n993), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1013), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1000), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1008), .B1(new_n1011), .B2(new_n1026), .ZN(new_n1027));
  AND4_X1   g602(.A1(new_n759), .A2(new_n1021), .A3(new_n1013), .A4(new_n1024), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n497), .B2(new_n993), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n947), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT45), .B(new_n993), .C1(new_n996), .C2(new_n997), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT111), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n497), .A2(new_n1034), .A3(KEYINPUT45), .A4(new_n993), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1013), .B(KEYINPUT110), .C1(new_n1017), .C2(KEYINPUT45), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1028), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1000), .B1(new_n1040), .B2(G168), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G168), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT63), .B1(new_n1027), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1011), .A2(new_n1026), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1011), .B2(new_n1026), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1025), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n947), .B1(new_n998), .B2(new_n945), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1048), .B2(new_n1014), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT109), .A3(new_n1010), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1046), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1044), .B1(new_n1042), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1008), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1002), .A2(new_n1003), .A3(new_n688), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1001), .B1(new_n1056), .B2(new_n981), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1043), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1046), .A2(new_n1051), .A3(new_n1044), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1008), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1028), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G286), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1041), .A3(KEYINPUT51), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  AOI211_X1 g642(.A(G286), .B(new_n1028), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n1000), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1065), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1031), .A2(new_n1036), .A3(new_n1037), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1018), .B2(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1021), .A2(new_n1013), .A3(new_n1024), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT121), .B(G1961), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1061), .A2(G168), .A3(new_n1062), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1040), .A2(G168), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1041), .A2(KEYINPUT51), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT120), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1065), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1091), .B2(KEYINPUT62), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1058), .B1(new_n1074), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1079), .A2(new_n748), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n999), .A2(new_n950), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT117), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1079), .A2(new_n748), .B1(new_n950), .B2(new_n999), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n603), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT117), .B(new_n602), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT113), .B1(G299), .B2(KEYINPUT112), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(G299), .B2(KEYINPUT113), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT113), .B(new_n1109), .C1(G299), .C2(KEYINPUT112), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1079), .A2(new_n744), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1018), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1018), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1119), .A2(new_n1115), .B1(new_n1079), .B2(new_n744), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G299), .A2(KEYINPUT112), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT57), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT61), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n998), .B2(new_n947), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1018), .B2(G1996), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(new_n1132), .C1(new_n1018), .C2(G1996), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n552), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1134), .A2(new_n1139), .A3(new_n552), .A4(new_n1136), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1126), .A2(new_n1130), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1107), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OR3_X1    g718(.A1(new_n1099), .A2(KEYINPUT114), .A3(new_n602), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT114), .B1(new_n1099), .B2(new_n602), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1127), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1146), .A2(KEYINPUT115), .A3(new_n1129), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT115), .B1(new_n1146), .B2(new_n1129), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1143), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1013), .A2(KEYINPUT122), .ZN(new_n1152));
  AND3_X1   g727(.A1(G160), .A2(KEYINPUT122), .A3(G40), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(new_n946), .A3(new_n1014), .A4(new_n1076), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT54), .B1(new_n1157), .B2(new_n1083), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1155), .A2(new_n1078), .A3(KEYINPUT123), .A4(new_n1081), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(G171), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1077), .A2(G301), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1163), .A2(KEYINPUT54), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n1059), .A3(new_n1008), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1158), .B(new_n1166), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1143), .A2(new_n1149), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1151), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1093), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n967), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n593), .B(G1986), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n949), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n972), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g751(.A(KEYINPUT124), .B(new_n1174), .C1(new_n1093), .C2(new_n1170), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n971), .B1(new_n1176), .B2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n1180));
  NOR2_X1   g754(.A1(G229), .A2(new_n460), .ZN(new_n1181));
  NOR2_X1   g755(.A1(G401), .A2(G227), .ZN(new_n1182));
  AND2_X1   g756(.A1(new_n860), .A2(new_n1182), .ZN(new_n1183));
  AND4_X1   g757(.A1(new_n1180), .A2(new_n940), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g758(.A(new_n1181), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1185), .B1(new_n938), .B2(new_n939), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1180), .B1(new_n1186), .B2(new_n1183), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1184), .A2(new_n1187), .ZN(G308));
  NAND3_X1  g762(.A1(new_n940), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n1186), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1191), .ZN(G225));
endmodule


