//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971;
  XNOR2_X1  g000(.A(G57gat), .B(G85gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G29gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT78), .B(G1gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G225gat), .A2(G233gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n212));
  OAI21_X1  g011(.A(G148gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G148gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n214), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n217), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G155gat), .B(G162gat), .Z(new_n226));
  AOI22_X1  g025(.A1(new_n215), .A2(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G113gat), .ZN(new_n233));
  INV_X1    g032(.A(G113gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237));
  INV_X1    g036(.A(G134gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G127gat), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n231), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n231), .B2(new_n239), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n227), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n228), .B1(new_n236), .B2(new_n237), .ZN(new_n245));
  AOI211_X1 g044(.A(KEYINPUT1), .B(G134gat), .C1(new_n233), .C2(new_n235), .ZN(new_n246));
  OAI21_X1  g045(.A(G127gat), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n239), .A3(new_n240), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(new_n227), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n210), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(new_n227), .C1(new_n241), .C2(new_n242), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT76), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n249), .B2(new_n227), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n209), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n243), .A2(new_n257), .A3(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n225), .A2(new_n226), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n211), .A2(new_n212), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n222), .B1(new_n260), .B2(G148gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n221), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n241), .A2(new_n242), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n227), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT5), .B(new_n251), .C1(new_n256), .C2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n271));
  INV_X1    g070(.A(new_n253), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n268), .B(new_n271), .C1(new_n272), .C2(new_n255), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n208), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n270), .A2(new_n208), .A3(new_n273), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(new_n275), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT80), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n207), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n270), .A2(new_n208), .A3(new_n273), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n276), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT25), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(KEYINPUT23), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n295), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n290), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n294), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(G176gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n297), .A2(KEYINPUT64), .ZN(new_n312));
  OAI211_X1 g111(.A(KEYINPUT23), .B(new_n296), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n303), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n304), .B1(new_n305), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n298), .A2(KEYINPUT26), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n301), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT27), .B(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT28), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT28), .B(new_n322), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n320), .B(new_n292), .C1(new_n323), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n330), .B(KEYINPUT72), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n321), .A2(new_n322), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n326), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(KEYINPUT66), .A3(new_n320), .A4(new_n292), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n305), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  INV_X1    g142(.A(new_n304), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n331), .A2(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n333), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT69), .B(G197gat), .ZN(new_n350));
  INV_X1    g149(.A(G204gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT70), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n355), .B(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n358), .B(new_n357), .C1(new_n352), .C2(new_n353), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n331), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n342), .A2(new_n344), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n368), .B2(new_n328), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT73), .B1(new_n369), .B2(new_n331), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n316), .B2(new_n329), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT73), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n332), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n366), .B1(new_n365), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G64gat), .ZN(new_n378));
  INV_X1    g177(.A(G92gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n288), .B(new_n289), .C1(new_n376), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(new_n346), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n316), .A2(new_n343), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n332), .B1(new_n385), .B2(new_n341), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n365), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n347), .A2(new_n348), .ZN(new_n388));
  INV_X1    g187(.A(new_n333), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n364), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n380), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT30), .B1(new_n392), .B2(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n380), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n381), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n287), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n362), .A2(new_n371), .A3(new_n363), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n266), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n263), .ZN(new_n400));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n401), .B(G22gat), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n227), .B2(new_n266), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n400), .B(new_n403), .C1(new_n365), .C2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n365), .A2(new_n404), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n227), .B1(new_n398), .B2(new_n266), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G50gat), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n405), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n405), .B2(new_n408), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n347), .A2(new_n249), .ZN(new_n416));
  INV_X1    g215(.A(G227gat), .ZN(new_n417));
  INV_X1    g216(.A(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n341), .B(new_n265), .C1(new_n345), .C2(new_n346), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n421), .B(KEYINPUT32), .C1(new_n423), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT34), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n420), .ZN(new_n433));
  INV_X1    g232(.A(new_n419), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT34), .B(new_n419), .C1(new_n416), .C2(new_n420), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT68), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n428), .A3(new_n430), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  INV_X1    g242(.A(new_n435), .ZN(new_n444));
  INV_X1    g243(.A(new_n436), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n428), .A2(new_n430), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT68), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n439), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n397), .A2(new_n415), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n372), .A2(new_n373), .A3(new_n332), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n373), .B1(new_n372), .B2(new_n332), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n364), .B1(new_n454), .B2(new_n367), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n455), .B2(new_n366), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n349), .A2(new_n365), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(KEYINPUT37), .C1(new_n375), .C2(new_n365), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n380), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT82), .ZN(new_n461));
  INV_X1    g260(.A(new_n380), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n387), .A2(new_n391), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n451), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n457), .A4(new_n459), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n376), .A2(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n457), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n392), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n284), .A2(new_n276), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n413), .A2(new_n414), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n268), .B1(new_n272), .B2(new_n255), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n210), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n244), .A2(new_n250), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n476), .B(KEYINPUT39), .C1(new_n210), .C2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(new_n208), .C1(KEYINPUT39), .C2(new_n476), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT40), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n395), .A2(new_n480), .A3(new_n282), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n437), .A2(new_n428), .A3(new_n430), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n483), .A2(new_n446), .A3(new_n415), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n287), .A2(new_n396), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n415), .B1(new_n442), .B2(new_n447), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n284), .A2(new_n276), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n395), .A2(new_n488), .A3(KEYINPUT35), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n450), .A2(new_n482), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT16), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(G1gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(G1gat), .B2(new_n492), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(G8gat), .Z(new_n496));
  XOR2_X1   g295(.A(G57gat), .B(G64gat), .Z(new_n497));
  AOI21_X1  g296(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G78gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(KEYINPUT89), .B2(new_n498), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505));
  NAND2_X1  g304(.A1(new_n497), .A2(KEYINPUT9), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n501), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT19), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT19), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G127gat), .B(G155gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(KEYINPUT91), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n510), .A2(KEYINPUT20), .A3(new_n512), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n522));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G183gat), .B(G211gat), .Z(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n525), .B(new_n526), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n518), .B1(new_n515), .B2(new_n519), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n521), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT84), .B(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  OR3_X1    g334(.A1(new_n534), .A2(KEYINPUT87), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT87), .B1(new_n534), .B2(new_n535), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT85), .B(G50gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(G43gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT86), .ZN(new_n542));
  NOR2_X1   g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545));
  OR2_X1    g344(.A1(G43gat), .A2(G50gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G43gat), .A2(G50gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n550), .B(new_n539), .C1(new_n540), .C2(G43gat), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n538), .A2(new_n542), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n534), .A2(new_n535), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n553), .B2(new_n544), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(KEYINPUT17), .A3(new_n554), .ZN(new_n558));
  XNOR2_X1  g357(.A(G99gat), .B(G106gat), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n379), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(new_n561), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n566), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT92), .A3(new_n559), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n557), .A2(new_n558), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n570), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n572), .A2(new_n576), .A3(new_n573), .A4(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(KEYINPUT93), .A3(new_n579), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n580), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n533), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT96), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n571), .A2(KEYINPUT94), .A3(new_n507), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n507), .A2(KEYINPUT94), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n506), .A2(new_n505), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n500), .B2(new_n503), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n600), .A3(new_n570), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT10), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n570), .A2(KEYINPUT10), .A3(new_n507), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT95), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n570), .A2(new_n605), .A3(KEYINPUT10), .A4(new_n507), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n594), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n595), .A2(new_n601), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT97), .A3(new_n593), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n601), .A3(new_n593), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n297), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n351), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n608), .A2(new_n610), .A3(new_n619), .A4(new_n613), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT98), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(KEYINPUT98), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n491), .A2(new_n591), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n557), .A2(new_n496), .A3(new_n558), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n495), .B(G8gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n555), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n626), .A2(KEYINPUT18), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n628), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n555), .A2(new_n627), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT18), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT88), .ZN(new_n641));
  XNOR2_X1  g440(.A(G169gat), .B(G197gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G113gat), .B(G141gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n637), .B(new_n640), .C1(new_n641), .C2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n641), .A3(new_n635), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  INV_X1    g449(.A(new_n640), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n636), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n625), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n287), .B(KEYINPUT99), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT100), .B(G1gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1324gat));
  AND2_X1   g457(.A1(new_n625), .A2(new_n653), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(KEYINPUT101), .A3(new_n395), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n654), .B2(new_n396), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n660), .B(new_n662), .C1(new_n663), .C2(G8gat), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n654), .B2(new_n396), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(KEYINPUT103), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(G1325gat));
  NAND2_X1  g473(.A1(new_n448), .A2(new_n449), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n659), .A2(G15gat), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n442), .A2(new_n447), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n659), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n654), .A2(new_n474), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n397), .A2(new_n415), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n482), .A2(new_n684), .A3(new_n675), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n278), .A2(KEYINPUT80), .A3(new_n279), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n284), .A2(new_n285), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n686), .A2(new_n687), .B1(new_n274), .B2(new_n275), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n439), .A2(new_n474), .A3(new_n441), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n688), .A2(new_n689), .A3(new_n395), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT35), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n490), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n590), .B1(new_n685), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n533), .A2(new_n624), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n693), .A2(new_n653), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n655), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n534), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT44), .B1(new_n491), .B2(new_n590), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n685), .A2(new_n692), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  INV_X1    g500(.A(new_n590), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n653), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n648), .A2(new_n652), .A3(KEYINPUT104), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n704), .A2(new_n694), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n655), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n698), .B1(new_n534), .B2(new_n711), .ZN(G1328gat));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n535), .A3(new_n395), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT46), .Z(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n710), .B2(new_n396), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n704), .A2(new_n676), .A3(new_n694), .A4(new_n709), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT47), .B1(new_n718), .B2(KEYINPUT105), .ZN(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n695), .A2(new_n720), .A3(new_n678), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n719), .B(new_n722), .ZN(G1330gat));
  INV_X1    g522(.A(new_n540), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n695), .A2(new_n724), .A3(new_n415), .ZN(new_n725));
  INV_X1    g524(.A(new_n710), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n415), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(new_n540), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT48), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n724), .B1(new_n726), .B2(new_n415), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n725), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1331gat));
  INV_X1    g532(.A(new_n624), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n491), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n709), .A2(new_n591), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n696), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n396), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n678), .B(KEYINPUT106), .Z(new_n747));
  NAND3_X1  g546(.A1(new_n738), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G71gat), .B1(new_n737), .B2(new_n675), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g550(.A1(new_n738), .A2(new_n415), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g552(.A1(new_n530), .A2(new_n532), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n708), .A2(KEYINPUT107), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n708), .B2(new_n754), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n693), .A2(KEYINPUT51), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT51), .B1(new_n693), .B2(new_n759), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n565), .A3(new_n696), .A4(new_n624), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n624), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n701), .B1(new_n700), .B2(new_n702), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT44), .B(new_n590), .C1(new_n685), .C2(new_n692), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT108), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n764), .B1(new_n699), .B2(new_n703), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n655), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n763), .B1(new_n773), .B2(new_n565), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT109), .B(new_n763), .C1(new_n773), .C2(new_n565), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1336gat));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n395), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(new_n779), .B2(G92gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n734), .A2(new_n396), .A3(G92gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n780), .A2(KEYINPUT111), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT111), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n760), .A2(new_n761), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n781), .B(KEYINPUT110), .Z(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n771), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT108), .B(new_n764), .C1(new_n699), .C2(new_n703), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n395), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n787), .B1(new_n790), .B2(G92gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n783), .A2(new_n784), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  AOI21_X1  g592(.A(new_n675), .B1(new_n769), .B2(new_n772), .ZN(new_n794));
  INV_X1    g593(.A(G99gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n678), .A2(new_n795), .A3(new_n624), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT112), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n795), .B1(new_n785), .B2(new_n797), .ZN(G1338gat));
  OAI21_X1  g597(.A(G106gat), .B1(new_n768), .B2(new_n474), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n734), .A2(G106gat), .A3(new_n474), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n799), .B(new_n800), .C1(new_n785), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(KEYINPUT113), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n760), .B2(new_n761), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT114), .B(new_n803), .C1(new_n760), .C2(new_n761), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n415), .B1(new_n788), .B2(new_n789), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(G106gat), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n802), .B1(new_n810), .B2(new_n800), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  INV_X1    g611(.A(new_n607), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n593), .C1(KEYINPUT10), .C2(new_n609), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n608), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n617), .B1(new_n608), .B2(KEYINPUT54), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n608), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n608), .A2(KEYINPUT54), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT55), .A4(new_n617), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n817), .A2(new_n620), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n706), .A3(new_n707), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n637), .A2(new_n647), .A3(new_n640), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n629), .B1(new_n626), .B2(new_n628), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n633), .A2(new_n634), .A3(new_n632), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n646), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(KEYINPUT115), .B(new_n646), .C1(new_n824), .C2(new_n825), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n823), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n623), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n621), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n702), .B1(new_n822), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n702), .A2(new_n821), .A3(new_n830), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n754), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n736), .A2(new_n734), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n655), .B(new_n395), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n487), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT116), .ZN(new_n839));
  INV_X1    g638(.A(new_n653), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n484), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n708), .A2(G113gat), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT117), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(G1340gat));
  OAI21_X1  g644(.A(G120gat), .B1(new_n839), .B2(new_n734), .ZN(new_n846));
  INV_X1    g645(.A(new_n842), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n232), .A3(new_n624), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1341gat));
  XNOR2_X1  g648(.A(KEYINPUT67), .B(G127gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n839), .B2(new_n754), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n754), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n842), .B2(new_n852), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n839), .B2(new_n590), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n238), .A3(new_n702), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  AOI21_X1  g657(.A(new_n474), .B1(new_n835), .B2(new_n836), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n655), .A2(new_n676), .A3(new_n395), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n840), .A2(G141gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n861), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n260), .ZN(new_n870));
  XNOR2_X1  g669(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n859), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n653), .A2(new_n620), .A3(new_n820), .A4(new_n817), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n702), .B1(new_n832), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n754), .B1(new_n875), .B2(new_n834), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n873), .B(new_n474), .C1(new_n836), .C2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n860), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n870), .B1(new_n878), .B2(new_n840), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n867), .A2(new_n868), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n869), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n709), .B(new_n860), .C1(new_n872), .C2(new_n877), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(new_n870), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n883), .B2(new_n870), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(new_n867), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(new_n880), .ZN(G1344gat));
  INV_X1    g687(.A(new_n861), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n223), .A3(new_n624), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n878), .B2(new_n734), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n223), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n702), .A2(new_n821), .A3(new_n830), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n821), .A2(new_n653), .B1(new_n624), .B2(new_n830), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n702), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n591), .A2(new_n624), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n896), .A2(new_n754), .B1(new_n840), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT122), .B(new_n873), .C1(new_n898), .C2(new_n474), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n840), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n474), .B1(new_n876), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n835), .A2(new_n836), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n415), .A3(new_n871), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n899), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n624), .A3(new_n860), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n891), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n890), .B1(new_n893), .B2(new_n908), .ZN(G1345gat));
  NOR3_X1   g708(.A1(new_n878), .A2(new_n219), .A3(new_n754), .ZN(new_n910));
  AOI21_X1  g709(.A(G155gat), .B1(new_n889), .B2(new_n533), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1346gat));
  NOR3_X1   g711(.A1(new_n878), .A2(new_n220), .A3(new_n590), .ZN(new_n913));
  AOI21_X1  g712(.A(G162gat), .B1(new_n889), .B2(new_n702), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  NAND3_X1  g714(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n655), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n696), .B1(new_n835), .B2(new_n836), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(KEYINPUT123), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n395), .B(new_n484), .C1(new_n917), .C2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n296), .B(new_n709), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n696), .A2(new_n396), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n904), .A2(new_n474), .A3(new_n747), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G169gat), .B1(new_n926), .B2(new_n840), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n928), .ZN(G1348gat));
  NOR4_X1   g728(.A1(new_n926), .A2(new_n311), .A3(new_n312), .A4(new_n734), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n624), .B1(new_n922), .B2(new_n923), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n297), .ZN(G1349gat));
  INV_X1    g731(.A(new_n321), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n920), .A2(new_n933), .A3(new_n754), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n926), .A2(new_n754), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G183gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n934), .A2(new_n937), .A3(KEYINPUT60), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT60), .B1(new_n934), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1350gat));
  OAI211_X1 g739(.A(new_n322), .B(new_n702), .C1(new_n922), .C2(new_n923), .ZN(new_n941));
  OAI21_X1  g740(.A(G190gat), .B1(new_n926), .B2(new_n590), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1351gat));
  OR2_X1    g743(.A1(new_n918), .A2(KEYINPUT123), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n396), .B1(new_n945), .B2(new_n916), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n676), .A2(new_n474), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n709), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n696), .A2(new_n676), .A3(new_n396), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n906), .A2(new_n653), .A3(new_n951), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n948), .A2(new_n950), .B1(new_n952), .B2(new_n949), .ZN(G1352gat));
  NAND4_X1  g752(.A1(new_n946), .A2(new_n351), .A3(new_n624), .A4(new_n947), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n906), .A2(new_n624), .A3(new_n951), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n955), .B(new_n956), .C1(new_n351), .C2(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n906), .A2(new_n533), .A3(new_n951), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G211gat), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT63), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(KEYINPUT126), .A3(new_n963), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n948), .A2(G211gat), .A3(new_n754), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n960), .A2(new_n966), .A3(new_n961), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(G1354gat));
  AND4_X1   g767(.A1(G218gat), .A2(new_n906), .A3(new_n702), .A4(new_n951), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n946), .A2(new_n702), .A3(new_n947), .ZN(new_n970));
  INV_X1    g769(.A(G218gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G1355gat));
endmodule


