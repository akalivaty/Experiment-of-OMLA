//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n642, new_n644, new_n645, new_n646, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1185,
    new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G137), .A4(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n462), .A2(KEYINPUT67), .A3(G137), .A4(new_n461), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G101), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT68), .B1(new_n466), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n461), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(G2104), .B2(new_n461), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n466), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G101), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n474), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n474), .A2(new_n485), .A3(KEYINPUT70), .A4(new_n481), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n465), .B1(new_n488), .B2(new_n489), .ZN(G160));
  NAND2_X1  g065(.A1(new_n467), .A2(new_n469), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n462), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(new_n461), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G136), .ZN(new_n497));
  OR2_X1    g072(.A1(G100), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n492), .A2(new_n494), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(new_n461), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(G124), .B2(new_n502), .ZN(G162));
  NAND4_X1  g078(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n462), .A2(G138), .A3(new_n461), .A4(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n509), .B1(KEYINPUT74), .B2(KEYINPUT4), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  AND2_X1   g086(.A1(G126), .A2(G2105), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n511), .B1(new_n462), .B2(new_n512), .ZN(new_n513));
  AND4_X1   g088(.A1(new_n511), .A2(new_n467), .A3(new_n469), .A4(new_n512), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n461), .A2(G114), .ZN(new_n515));
  OAI21_X1  g090(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n461), .A2(G114), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n519), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n513), .A2(new_n514), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n510), .A2(new_n522), .ZN(G164));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(G62), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(new_n527), .ZN(new_n532));
  INV_X1    g107(.A(G62), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT76), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT75), .B(G651), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT75), .B(G651), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT6), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n528), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G88), .ZN(new_n543));
  INV_X1    g118(.A(G50), .ZN(new_n544));
  OAI211_X1 g119(.A(G543), .B(new_n541), .C1(new_n536), .C2(new_n540), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n537), .A2(new_n546), .ZN(G166));
  INV_X1    g122(.A(new_n545), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G51), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  INV_X1    g127(.A(G89), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n549), .B(new_n550), .C1(new_n556), .C2(new_n557), .ZN(G286));
  INV_X1    g133(.A(G286), .ZN(G168));
  INV_X1    g134(.A(new_n542), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G90), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n548), .A2(G52), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n538), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(G301));
  INV_X1    g140(.A(G301), .ZN(G171));
  NAND2_X1  g141(.A1(new_n560), .A2(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n548), .A2(G43), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n538), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  AND3_X1   g148(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G36), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G188));
  NAND4_X1  g153(.A1(new_n539), .A2(G53), .A3(G543), .A4(new_n541), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT79), .B1(new_n579), .B2(KEYINPUT9), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  INV_X1    g156(.A(G53), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n545), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n586), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n579), .A2(KEYINPUT78), .A3(KEYINPUT9), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n580), .A2(new_n585), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G78), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G65), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n532), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G91), .B2(new_n560), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n589), .A2(new_n595), .ZN(G299));
  INV_X1    g171(.A(G166), .ZN(G303));
  NAND4_X1  g172(.A1(new_n539), .A2(G87), .A3(new_n528), .A4(new_n541), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G49), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT81), .B1(new_n545), .B2(new_n601), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n545), .A2(KEYINPUT81), .A3(new_n601), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT82), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n600), .A2(new_n606), .A3(new_n602), .A4(new_n603), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G288));
  NAND3_X1  g183(.A1(new_n548), .A2(KEYINPUT84), .A3(G48), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n528), .A2(G61), .ZN(new_n610));
  NAND2_X1  g185(.A1(G73), .A2(G543), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT83), .Z(new_n612));
  OAI21_X1  g187(.A(new_n536), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n539), .A2(G86), .A3(new_n528), .A4(new_n541), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n615));
  INV_X1    g190(.A(G48), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n545), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n609), .A2(new_n613), .A3(new_n614), .A4(new_n617), .ZN(G305));
  INV_X1    g193(.A(G85), .ZN(new_n619));
  INV_X1    g194(.A(G47), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n542), .A2(new_n619), .B1(new_n620), .B2(new_n545), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(new_n538), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(G301), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  OR3_X1    g203(.A1(new_n542), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(G79), .A2(G543), .ZN(new_n630));
  INV_X1    g205(.A(G66), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n532), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n548), .A2(G54), .B1(G651), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT10), .B1(new_n542), .B2(new_n628), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n629), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n627), .B1(new_n635), .B2(G868), .ZN(G284));
  OAI21_X1  g211(.A(new_n627), .B1(new_n635), .B2(G868), .ZN(G321));
  NAND2_X1  g212(.A1(G286), .A2(G868), .ZN(new_n638));
  INV_X1    g213(.A(G299), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(G868), .B2(new_n639), .ZN(G297));
  OAI21_X1  g215(.A(new_n638), .B1(G868), .B2(new_n639), .ZN(G280));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n635), .B1(new_n642), .B2(G860), .ZN(G148));
  NOR2_X1   g218(.A1(new_n572), .A2(G868), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G868), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(G323));
  XNOR2_X1  g222(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n648));
  XNOR2_X1  g223(.A(G323), .B(new_n648), .ZN(G282));
  NAND2_X1  g224(.A1(new_n502), .A2(G123), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n496), .A2(G135), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(KEYINPUT89), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(KEYINPUT89), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n653), .B(new_n654), .C1(G111), .C2(new_n461), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G2096), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(KEYINPUT88), .B2(G2100), .ZN(new_n658));
  NAND2_X1  g233(.A1(KEYINPUT88), .A2(G2100), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n476), .A2(new_n478), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(new_n462), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT12), .Z(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT13), .Z(new_n663));
  AOI21_X1  g238(.A(new_n658), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  OAI221_X1 g239(.A(new_n664), .B1(G2096), .B2(new_n656), .C1(new_n659), .C2(new_n663), .ZN(G156));
  XNOR2_X1  g240(.A(G2427), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2430), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT15), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(G2435), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(G2435), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(KEYINPUT14), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2443), .B(G2446), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1341), .B(G1348), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2451), .B(G2454), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G14), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G401));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT91), .B(KEYINPUT17), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2067), .B(G2678), .Z(new_n685));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n689), .A2(new_n686), .ZN(new_n690));
  INV_X1    g265(.A(new_n685), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n682), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n682), .A2(new_n691), .A3(new_n686), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT18), .Z(new_n694));
  NAND3_X1  g269(.A1(new_n688), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  XNOR2_X1  g271(.A(G2096), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT19), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n709), .B(new_n710), .C1(new_n708), .C2(new_n707), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n711), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1991), .B(G1996), .ZN(new_n716));
  INV_X1    g291(.A(G1981), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n715), .B(new_n719), .ZN(G229));
  NOR2_X1   g295(.A1(G6), .A2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G305), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT96), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G23), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n726), .A2(G16), .A3(G23), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n727), .B(new_n728), .C1(new_n604), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n729), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n725), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT34), .Z(new_n739));
  INV_X1    g314(.A(G290), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G16), .B2(G24), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(new_n713), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n713), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(G25), .ZN(new_n746));
  INV_X1    g321(.A(new_n502), .ZN(new_n747));
  INV_X1    g322(.A(G119), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n747), .A2(KEYINPUT95), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n461), .A2(G107), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n496), .A2(G131), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT95), .B1(new_n747), .B2(new_n748), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT35), .B(G1991), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n756), .B(new_n757), .Z(new_n758));
  NOR3_X1   g333(.A1(new_n743), .A2(new_n744), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n739), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT36), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n729), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n635), .B2(new_n729), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT98), .B(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n763), .B(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G19), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n572), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT100), .B(G1341), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n745), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n745), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G168), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G16), .B2(G21), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n656), .A2(new_n745), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(KEYINPUT103), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G35), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G162), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT29), .B(G2090), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT31), .B(G11), .Z(new_n786));
  NOR3_X1   g361(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AND4_X1   g362(.A1(new_n774), .A2(new_n778), .A3(new_n780), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n776), .A2(new_n777), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT104), .ZN(new_n790));
  OR2_X1    g365(.A1(KEYINPUT24), .A2(G34), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT24), .A2(G34), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n791), .A2(new_n745), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G160), .B2(new_n745), .ZN(new_n794));
  INV_X1    g369(.A(G2084), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G28), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(G28), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n798), .A2(new_n799), .A3(new_n745), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n788), .A2(new_n790), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(G171), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G5), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT105), .Z(new_n806));
  NAND3_X1  g381(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT25), .Z(new_n808));
  INV_X1    g383(.A(G139), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n495), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT101), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(KEYINPUT101), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n811), .A2(new_n812), .B1(new_n461), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT102), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G29), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G29), .B2(G33), .ZN(new_n817));
  INV_X1    g392(.A(G2072), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n803), .A2(new_n804), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n745), .A2(G26), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n502), .A2(G128), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n496), .A2(G140), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n461), .A2(G116), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n821), .B1(new_n826), .B2(G29), .ZN(new_n827));
  MUX2_X1   g402(.A(new_n821), .B(new_n827), .S(KEYINPUT28), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2067), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n806), .A2(new_n819), .A3(new_n820), .A4(new_n829), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n729), .A2(KEYINPUT23), .A3(G20), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT23), .B1(new_n729), .B2(G20), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n831), .B(new_n832), .C1(G299), .C2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1956), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n834), .B1(KEYINPUT103), .B2(new_n779), .C1(new_n817), .C2(new_n818), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n801), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n761), .A2(new_n766), .A3(new_n770), .A4(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT106), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n502), .A2(G129), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n496), .A2(G141), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n660), .A2(G105), .ZN(new_n841));
  NAND3_X1  g416(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT26), .Z(new_n843));
  NAND4_X1  g418(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  MUX2_X1   g419(.A(G32), .B(new_n844), .S(G29), .Z(new_n845));
  XOR2_X1   g420(.A(KEYINPUT27), .B(G1996), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OR3_X1    g422(.A1(new_n837), .A2(new_n838), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n838), .B1(new_n837), .B2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G311));
  OR2_X1    g425(.A1(new_n837), .A2(new_n847), .ZN(G150));
  AOI22_X1  g426(.A1(new_n560), .A2(G93), .B1(G55), .B2(new_n548), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT107), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n854), .B2(new_n538), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n571), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n572), .A2(new_n855), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n635), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n857), .B1(new_n865), .B2(G860), .ZN(G145));
  XNOR2_X1  g441(.A(new_n755), .B(new_n656), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n815), .A2(new_n826), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n815), .A2(new_n826), .ZN(new_n870));
  XNOR2_X1  g445(.A(G164), .B(new_n662), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n815), .A2(new_n826), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n871), .B1(new_n874), .B2(new_n868), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n867), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n872), .B1(new_n869), .B2(new_n870), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n868), .A3(new_n871), .ZN(new_n878));
  INV_X1    g453(.A(new_n867), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(G162), .B(G160), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n502), .A2(G130), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n496), .A2(G142), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(KEYINPUT108), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(KEYINPUT108), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n886), .B(new_n887), .C1(G118), .C2(new_n461), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n844), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n882), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n876), .A2(new_n891), .A3(new_n880), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT109), .B(G37), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g473(.A1(new_n858), .A2(G868), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n861), .B(new_n645), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n635), .B1(G299), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n901), .B2(G299), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n639), .A2(KEYINPUT110), .A3(new_n635), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT41), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n909), .B2(new_n900), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(G303), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n623), .A2(G166), .A3(new_n625), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n604), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n604), .A3(new_n913), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n916), .A2(new_n722), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n722), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n910), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n899), .B1(new_n926), .B2(G868), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT111), .ZN(G295));
  NAND2_X1  g503(.A1(new_n926), .A2(G868), .ZN(new_n929));
  INV_X1    g504(.A(new_n899), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n905), .A2(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n907), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(G286), .A2(G171), .ZN(new_n936));
  NOR2_X1   g511(.A1(G286), .A2(G171), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n861), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n556), .A2(new_n557), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(new_n549), .A3(new_n550), .A4(G301), .ZN(new_n943));
  NAND2_X1  g518(.A1(G286), .A2(G171), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n860), .A3(new_n859), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n938), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n933), .B(new_n935), .C1(new_n941), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n938), .A2(new_n945), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(new_n907), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n920), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n895), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(KEYINPUT112), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n905), .A3(new_n940), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n933), .A2(new_n935), .A3(new_n948), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n920), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n940), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n949), .B1(new_n958), .B2(new_n908), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT113), .B1(new_n959), .B2(new_n920), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n932), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n955), .A2(new_n956), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n918), .B2(new_n919), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n966), .A3(new_n957), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n967), .B2(KEYINPUT43), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n967), .A2(new_n963), .A3(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n953), .A2(new_n971), .A3(new_n957), .A4(new_n960), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n932), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(new_n465), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n479), .B(KEYINPUT69), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT70), .B1(new_n978), .B2(new_n474), .ZN(new_n979));
  AND4_X1   g554(.A1(KEYINPUT70), .A2(new_n474), .A3(new_n481), .A4(new_n485), .ZN(new_n980));
  OAI211_X1 g555(.A(G40), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT115), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n983));
  NAND3_X1  g558(.A1(G160), .A2(new_n983), .A3(G40), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n510), .B2(new_n522), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n740), .A2(new_n713), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT116), .Z(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n713), .B2(new_n740), .ZN(new_n996));
  INV_X1    g571(.A(G2067), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n826), .B(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n844), .B(G1996), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n755), .A2(new_n757), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n755), .A2(new_n757), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n992), .B1(new_n996), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n986), .C1(new_n510), .C2(new_n522), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT117), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n987), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n981), .A2(KEYINPUT115), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n983), .B1(G160), .B2(G40), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G2090), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n986), .C1(new_n510), .C2(new_n522), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n989), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n982), .B2(new_n984), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G1971), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1010), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n985), .A2(new_n1014), .A3(new_n1012), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1027), .A2(G2090), .B1(G1971), .B2(new_n1023), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1010), .B1(new_n1028), .B2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n987), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n604), .A2(new_n1032), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1031), .A2(G8), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n613), .A2(new_n614), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(new_n717), .A3(new_n617), .A4(new_n609), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1031), .A3(G8), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n987), .B1(new_n982), .B2(new_n984), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1034), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1036), .B(new_n1043), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1026), .A2(new_n1029), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  AND3_X1   g626(.A1(G299), .A2(new_n1051), .A3(KEYINPUT57), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(KEYINPUT57), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(KEYINPUT57), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(G299), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1014), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n982), .B2(new_n984), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1956), .B1(new_n1059), .B2(new_n1012), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n1022), .B(new_n1062), .C1(new_n982), .C2(new_n984), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1057), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1023), .A2(new_n1061), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1012), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n1058), .C1(new_n982), .C2(new_n984), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1065), .B(new_n1066), .C1(new_n1068), .C2(G1956), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1064), .A2(KEYINPUT61), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT61), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1023), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT58), .B(G1341), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1073), .A2(G1996), .B1(new_n1044), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n572), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT59), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n997), .B(new_n1030), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n982), .B2(new_n984), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT60), .B(new_n1078), .C1(new_n1080), .C2(G1348), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT124), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(KEYINPUT124), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n635), .ZN(new_n1084));
  INV_X1    g659(.A(new_n635), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(KEYINPUT124), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1019), .A2(new_n1088), .B1(new_n1044), .B2(new_n997), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1072), .B(new_n1077), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1064), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1069), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1019), .B2(G2084), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1080), .A2(KEYINPUT121), .A3(new_n795), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1073), .A2(new_n777), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G286), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n1101), .B2(KEYINPUT125), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1102), .C1(new_n1099), .C2(G286), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(G8), .A3(G286), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1022), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n985), .A2(new_n773), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1019), .A2(new_n804), .ZN(new_n1112));
  OR4_X1    g687(.A1(new_n1110), .A2(new_n1022), .A3(new_n981), .A4(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1111), .A2(new_n1112), .A3(G301), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT126), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1110), .A2(new_n1109), .B1(new_n1019), .B2(new_n804), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(G301), .A4(new_n1113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1023), .A2(KEYINPUT53), .A3(new_n773), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1111), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G171), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1115), .A2(new_n1118), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(G301), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1116), .A2(G171), .A3(new_n1113), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(KEYINPUT54), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1107), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1094), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1107), .A2(KEYINPUT62), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1104), .A2(new_n1131), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1130), .A2(G171), .A3(new_n1120), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1050), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1099), .A2(G8), .A3(G168), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1029), .A2(new_n1048), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1025), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1048), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(G8), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1009), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1031), .A2(G8), .A3(new_n1035), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT52), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(KEYINPUT119), .A3(new_n1043), .A4(new_n1036), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1142), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1025), .A2(KEYINPUT63), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1136), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1139), .A2(new_n1140), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1142), .A2(new_n1026), .A3(new_n1147), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT120), .Z(new_n1154));
  OAI21_X1  g729(.A(new_n1038), .B1(new_n1154), .B2(new_n1042), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(G8), .A3(new_n1031), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1135), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1157), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n1049), .B2(new_n1137), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT122), .B(new_n1159), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1006), .B1(new_n1134), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n826), .A2(G2067), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n991), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  OR3_X1    g743(.A1(new_n991), .A2(new_n1168), .A3(G1996), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n992), .B1(new_n844), .B2(new_n999), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n991), .B2(G1996), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT47), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1005), .A2(new_n992), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n994), .A2(new_n992), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT48), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1167), .B(new_n1173), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1164), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G229), .ZN(new_n1180));
  AND2_X1   g754(.A1(new_n897), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g755(.A(G319), .ZN(new_n1182));
  NOR3_X1   g756(.A1(G401), .A2(new_n1182), .A3(G227), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n974), .A2(new_n1181), .A3(new_n1183), .ZN(G225));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1185));
  NAND2_X1  g759(.A1(G225), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g760(.A1(new_n974), .A2(new_n1181), .A3(new_n1183), .A4(KEYINPUT127), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1187), .ZN(G308));
endmodule


