//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  XNOR2_X1  g000(.A(KEYINPUT11), .B(G169gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G141gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT86), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n207), .A2(G43gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT15), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(G50gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n217), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT87), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT14), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n214), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n216), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n224), .B2(new_n220), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT17), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n230));
  INV_X1    g029(.A(new_n224), .ZN(new_n231));
  INV_X1    g030(.A(new_n213), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT86), .B(G50gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(new_n211), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n230), .B(new_n231), .C1(KEYINPUT15), .C2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n227), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G15gat), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G15gat), .A2(G22gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G1gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT88), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT88), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT16), .B1(new_n246), .B2(G1gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n241), .A2(new_n244), .A3(new_n242), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G8gat), .ZN(new_n252));
  INV_X1    g051(.A(G8gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n248), .A2(new_n249), .A3(new_n253), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G229gat), .A2(G233gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n227), .A2(new_n235), .B1(new_n252), .B2(new_n254), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT18), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n206), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n225), .A2(new_n228), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n258), .B(KEYINPUT13), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n259), .B1(new_n238), .B2(new_n256), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT18), .A3(new_n258), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n263), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n206), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT18), .B1(new_n272), .B2(new_n258), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(KEYINPUT90), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n255), .B1(new_n229), .B2(new_n237), .ZN(new_n279));
  INV_X1    g078(.A(new_n258), .ZN(new_n280));
  NOR4_X1   g079(.A1(new_n279), .A2(new_n262), .A3(new_n259), .A4(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n271), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G155gat), .B(G162gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(KEYINPUT2), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G141gat), .B(G148gat), .Z(new_n289));
  XNOR2_X1  g088(.A(G155gat), .B(G162gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT2), .B1(new_n291), .B2(KEYINPUT76), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT73), .B(G204gat), .Z(new_n296));
  INV_X1    g095(.A(G197gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT73), .B(G204gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G197gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G211gat), .B(G218gat), .Z(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n298), .A2(new_n308), .A3(new_n302), .A4(new_n304), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n307), .C2(new_n309), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n294), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(new_n309), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n288), .A2(new_n293), .A3(new_n295), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(KEYINPUT29), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n288), .A2(new_n293), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n315), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n240), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT31), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(new_n207), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT83), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n322), .A2(new_n326), .A3(new_n240), .A4(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G22gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n331), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT27), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT67), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT67), .B1(new_n344), .B2(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n341), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n343), .A2(new_n345), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT28), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(KEYINPUT26), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n353), .A2(new_n355), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G176gat), .ZN(new_n362));
  AND2_X1   g161(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT23), .B(new_n362), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT65), .B1(new_n356), .B2(KEYINPUT23), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n369), .B(new_n370), .C1(G169gat), .C2(G176gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n358), .A3(new_n371), .ZN(new_n372));
  OAI22_X1  g171(.A1(new_n367), .A2(new_n372), .B1(KEYINPUT66), .B2(new_n366), .ZN(new_n373));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n354), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT24), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT66), .B1(new_n376), .B2(new_n377), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n368), .A2(new_n358), .A3(new_n371), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n356), .A2(KEYINPUT23), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT25), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n361), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G113gat), .B(G120gat), .Z(new_n386));
  INV_X1    g185(.A(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT69), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(KEYINPUT1), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(KEYINPUT1), .ZN(new_n391));
  INV_X1    g190(.A(G127gat), .ZN(new_n392));
  INV_X1    g191(.A(G134gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G127gat), .A2(G134gat), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n390), .A2(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT68), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n388), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n394), .B(new_n395), .C1(new_n397), .C2(KEYINPUT1), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G227gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(KEYINPUT25), .A2(new_n383), .B1(new_n373), .B2(new_n378), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n399), .A2(new_n400), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n361), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n402), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT34), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n402), .A2(new_n409), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT70), .B1(new_n413), .B2(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n415));
  AOI211_X1 g214(.A(new_n415), .B(new_n406), .C1(new_n402), .C2(new_n409), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT32), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n414), .B2(new_n416), .ZN(new_n419));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  OAI221_X1 g223(.A(KEYINPUT32), .B1(new_n418), .B2(new_n424), .C1(new_n414), .C2(new_n416), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(KEYINPUT71), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT72), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n412), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n427), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n423), .A2(new_n425), .B1(KEYINPUT71), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n340), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT80), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n401), .A2(new_n294), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n399), .A2(new_n400), .B1(new_n288), .B2(new_n293), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT77), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n324), .A2(new_n400), .A3(new_n399), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n401), .A3(new_n319), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n438), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n401), .A2(new_n294), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n445), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT77), .A3(new_n439), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT78), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n455), .A2(KEYINPUT5), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n455), .B2(KEYINPUT5), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n437), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n458), .A2(new_n459), .A3(new_n437), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(new_n437), .C1(new_n458), .C2(new_n459), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n459), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n455), .A2(KEYINPUT5), .A3(new_n457), .ZN(new_n468));
  INV_X1    g267(.A(new_n437), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n385), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n407), .B2(new_n361), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n318), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n385), .A2(new_n474), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n472), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n473), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT75), .B1(new_n385), .B2(new_n473), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n480), .B(new_n317), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT74), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(new_n318), .C1(new_n475), .C2(new_n476), .ZN(new_n485));
  XOR2_X1   g284(.A(G8gat), .B(G36gat), .Z(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G64gat), .ZN(new_n487));
  INV_X1    g286(.A(G92gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n478), .A2(new_n483), .A3(new_n485), .A4(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n489), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n492), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n471), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT35), .B1(new_n431), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n412), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n423), .A2(new_n501), .A3(new_n425), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n423), .B2(new_n425), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n497), .B1(new_n466), .B2(new_n470), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n340), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n453), .A2(new_n439), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT84), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n439), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT39), .B(new_n512), .C1(new_n515), .C2(new_n511), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n439), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n516), .B(new_n437), .C1(KEYINPUT39), .C2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT40), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n497), .A3(new_n462), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT38), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n494), .A2(new_n521), .A3(new_n490), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n494), .A2(KEYINPUT37), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n478), .A2(new_n483), .A3(new_n485), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n490), .B1(new_n527), .B2(KEYINPUT38), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n480), .B(new_n318), .C1(new_n481), .C2(new_n482), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n317), .B1(new_n475), .B2(new_n476), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(KEYINPUT37), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n521), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n522), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n340), .B(new_n520), .C1(new_n533), .C2(new_n471), .ZN(new_n534));
  INV_X1    g333(.A(new_n340), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n499), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n504), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n502), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n426), .A2(new_n427), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n430), .B1(new_n540), .B2(new_n501), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(new_n536), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n285), .B1(new_n510), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G211gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT21), .ZN(new_n551));
  XOR2_X1   g350(.A(G57gat), .B(G64gat), .Z(new_n552));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553));
  INV_X1    g352(.A(G71gat), .ZN(new_n554));
  INV_X1    g353(.A(G78gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n558), .A3(new_n556), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n256), .B(new_n344), .C1(new_n551), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n551), .ZN(new_n564));
  OAI21_X1  g363(.A(G183gat), .B1(new_n564), .B2(new_n255), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n562), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n570), .ZN(new_n573));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT92), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n550), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n577), .A3(new_n549), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n586), .B2(new_n488), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n586), .B2(new_n488), .ZN(new_n589));
  NAND3_X1  g388(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n587), .A2(new_n592), .A3(new_n589), .A4(new_n590), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT93), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n597), .A3(new_n593), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n238), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n600), .B2(new_n266), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n584), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  INV_X1    g406(.A(new_n584), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n601), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n606), .A2(new_n609), .A3(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n583), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n596), .A2(new_n562), .A3(new_n598), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT94), .B(KEYINPUT10), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n560), .A2(new_n594), .A3(new_n561), .A4(new_n595), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n620), .A2(new_n625), .A3(new_n621), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n567), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n620), .B2(new_n622), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n362), .ZN(new_n636));
  INV_X1    g435(.A(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n640), .A3(new_n633), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n619), .A2(KEYINPUT97), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n617), .B1(new_n580), .B2(new_n582), .ZN(new_n645));
  INV_X1    g444(.A(new_n642), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n545), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n471), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g451(.A1(new_n545), .A2(new_n498), .A3(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n654));
  OR2_X1    g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n658), .B(new_n659), .C1(new_n253), .C2(new_n653), .ZN(G1325gat));
  AOI21_X1  g459(.A(G15gat), .B1(new_n649), .B2(new_n506), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n542), .A2(new_n239), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n649), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n649), .A2(new_n535), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n583), .A2(new_n642), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n617), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT98), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n544), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(G29gat), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n668), .A2(KEYINPUT98), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n650), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n534), .A2(new_n536), .A3(new_n542), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n507), .B(new_n340), .C1(new_n428), .C2(new_n430), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n340), .B(new_n508), .C1(new_n503), .C2(new_n504), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n678), .A2(KEYINPUT35), .B1(new_n507), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n617), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n618), .B1(new_n510), .B2(new_n543), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n284), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n275), .A2(new_n283), .A3(KEYINPUT100), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n667), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT101), .Z(new_n693));
  AND3_X1   g492(.A1(new_n684), .A2(new_n686), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(new_n650), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n675), .B(new_n676), .C1(new_n695), .C2(new_n671), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n697));
  INV_X1    g496(.A(G36gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n694), .B2(new_n497), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n544), .A2(new_n672), .A3(new_n669), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n497), .A2(new_n698), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n700), .A2(KEYINPUT46), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT46), .B1(new_n700), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n697), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n510), .A2(new_n543), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n706), .B2(new_n617), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n683), .B(new_n618), .C1(new_n510), .C2(new_n543), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n497), .A3(new_n693), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G36gat), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n711), .A2(KEYINPUT102), .A3(new_n703), .A4(new_n702), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n712), .ZN(G1329gat));
  NOR3_X1   g512(.A1(new_n700), .A2(G43gat), .A3(new_n505), .ZN(new_n714));
  INV_X1    g513(.A(new_n542), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n684), .A2(new_n715), .A3(new_n686), .A4(new_n693), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(G43gat), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g517(.A1(new_n684), .A2(new_n535), .A3(new_n686), .A4(new_n693), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n233), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n721));
  INV_X1    g520(.A(new_n233), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n544), .A2(new_n723), .A3(new_n672), .A4(new_n669), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n721), .A2(new_n535), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT105), .Z(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n720), .A2(new_n725), .A3(new_n729), .A4(new_n726), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n691), .A2(new_n619), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n706), .A2(new_n642), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n706), .A2(new_n737), .A3(new_n642), .A4(new_n734), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n650), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n736), .A2(new_n738), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n497), .B(KEYINPUT107), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  AOI21_X1  g548(.A(G71gat), .B1(new_n739), .B2(new_n506), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n715), .A2(G71gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT50), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n554), .B1(new_n742), .B2(new_n505), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n754), .B(new_n755), .C1(new_n742), .C2(new_n751), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(G1334gat));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n340), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT108), .B(G78gat), .Z(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n691), .A2(new_n583), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n684), .A2(new_n642), .A3(new_n686), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n471), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n471), .A2(G85gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n706), .A2(new_n617), .A3(new_n761), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n685), .B2(new_n761), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n642), .B(new_n764), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n763), .A2(new_n772), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n762), .B2(new_n744), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n744), .A2(G92gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n642), .B(new_n777), .C1(new_n767), .C2(new_n768), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  AOI211_X1 g578(.A(KEYINPUT110), .B(new_n766), .C1(new_n685), .C2(new_n761), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n765), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n782), .A3(new_n646), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n709), .A2(new_n497), .A3(new_n642), .A4(new_n761), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n783), .A2(new_n777), .B1(new_n784), .B2(G92gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n779), .B1(new_n785), .B2(new_n776), .ZN(G1337gat));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n762), .A2(new_n787), .A3(new_n542), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n762), .B2(new_n542), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(G99gat), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n765), .B(new_n766), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n505), .A2(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n642), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1338gat));
  NAND4_X1  g593(.A1(new_n709), .A2(new_n535), .A3(new_n642), .A4(new_n761), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n340), .A2(G106gat), .A3(new_n646), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT53), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n780), .A2(new_n782), .ZN(new_n800));
  AOI22_X1  g599(.A1(G106gat), .A2(new_n795), .B1(new_n800), .B2(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1339gat));
  INV_X1    g602(.A(new_n583), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  INV_X1    g604(.A(new_n628), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n624), .B2(new_n626), .ZN(new_n807));
  INV_X1    g606(.A(new_n630), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n631), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n627), .B2(new_n628), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n640), .B1(new_n811), .B2(new_n805), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT55), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n641), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n812), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n814), .A2(new_n688), .A3(new_n689), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n272), .A2(new_n258), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n268), .A2(new_n270), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n205), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n282), .A2(new_n206), .A3(new_n271), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n642), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n617), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n810), .B2(new_n812), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n274), .B2(new_n276), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n814), .A2(new_n827), .A3(new_n617), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n804), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n645), .A2(new_n690), .A3(KEYINPUT112), .A4(new_n646), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n645), .A2(new_n690), .A3(new_n646), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(new_n340), .A3(new_n506), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n743), .A2(new_n471), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n284), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT113), .B1(new_n837), .B2(G113gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n650), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n431), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n744), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n690), .A2(G113gat), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n838), .A2(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  NAND2_X1  g643(.A1(new_n835), .A2(new_n836), .ZN(new_n845));
  OAI21_X1  g644(.A(G120gat), .B1(new_n845), .B2(new_n646), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n842), .A2(G120gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n646), .ZN(G1341gat));
  NOR3_X1   g647(.A1(new_n845), .A2(new_n392), .A3(new_n804), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n841), .A2(new_n583), .A3(new_n744), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n392), .ZN(G1342gat));
  NOR2_X1   g650(.A1(new_n497), .A2(new_n618), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n841), .A2(new_n393), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n845), .B2(new_n618), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(G1343gat));
  AND2_X1   g659(.A1(new_n542), .A2(new_n535), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT115), .B1(new_n715), .B2(new_n340), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n863), .A2(new_n834), .A3(new_n864), .A4(new_n650), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(G141gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n284), .A4(new_n744), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n834), .A2(new_n869), .A3(new_n535), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n833), .A2(new_n830), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n817), .A2(new_n284), .A3(new_n641), .A4(new_n813), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n823), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n618), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n814), .A2(new_n827), .A3(new_n617), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n583), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n535), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT57), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n836), .A2(new_n542), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n870), .A2(new_n878), .A3(new_n691), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G141gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n868), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT116), .B1(new_n882), .B2(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n884), .B(new_n885), .C1(new_n868), .C2(new_n881), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n870), .A2(new_n878), .A3(new_n879), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n867), .B1(new_n887), .B2(new_n284), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n885), .ZN(new_n889));
  OAI22_X1  g688(.A1(new_n883), .A2(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n865), .A2(new_n743), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n642), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n617), .B1(new_n872), .B2(new_n823), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT117), .B1(new_n895), .B2(new_n828), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n826), .B1(new_n641), .B2(new_n639), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n816), .A2(new_n815), .B1(new_n275), .B2(new_n283), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n814), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n897), .B(new_n875), .C1(new_n900), .C2(new_n617), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n901), .A3(new_n804), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n285), .B1(new_n643), .B2(new_n647), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT118), .B(new_n869), .C1(new_n904), .C2(new_n340), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n834), .A2(KEYINPUT57), .A3(new_n535), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n340), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n642), .A3(new_n879), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n894), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT59), .B(new_n892), .C1(new_n887), .C2(new_n642), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n893), .B1(new_n912), .B2(new_n913), .ZN(G1345gat));
  AOI21_X1  g713(.A(G155gat), .B1(new_n891), .B2(new_n583), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n583), .A2(G155gat), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT119), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n887), .B2(new_n917), .ZN(G1346gat));
  XNOR2_X1  g717(.A(KEYINPUT76), .B(G162gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n866), .A2(new_n852), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n887), .A2(new_n617), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT120), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n919), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n650), .A2(new_n498), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n835), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n285), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT124), .B(G169gat), .C1(new_n925), .C2(new_n285), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n834), .A2(new_n471), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n834), .A2(KEYINPUT121), .A3(new_n471), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n744), .A2(new_n431), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT122), .Z(new_n938));
  AND2_X1   g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n363), .A2(new_n364), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n690), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n931), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n936), .A2(new_n938), .ZN(new_n943));
  INV_X1    g742(.A(new_n941), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n943), .A2(KEYINPUT123), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n930), .B1(new_n942), .B2(new_n945), .ZN(G1348gat));
  NOR3_X1   g745(.A1(new_n925), .A2(new_n362), .A3(new_n646), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n939), .A2(new_n642), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n362), .ZN(G1349gat));
  OAI21_X1  g748(.A(G183gat), .B1(new_n925), .B2(new_n804), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n583), .A2(new_n351), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n950), .B(new_n954), .C1(new_n943), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n925), .B2(new_n618), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(KEYINPUT125), .B(G190gat), .C1(new_n925), .C2(new_n618), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(KEYINPUT61), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n348), .A3(new_n617), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(G1351gat));
  NAND4_X1  g764(.A1(new_n934), .A2(new_n743), .A3(new_n861), .A4(new_n935), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(new_n297), .A3(new_n691), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n542), .A2(new_n924), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n910), .A2(new_n284), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n970), .B2(new_n297), .ZN(G1352gat));
  AND3_X1   g770(.A1(new_n934), .A2(new_n743), .A3(new_n935), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n972), .A2(new_n637), .A3(new_n861), .A4(new_n974), .ZN(new_n975));
  OAI22_X1  g774(.A1(new_n975), .A2(new_n646), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n966), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n977), .A2(new_n637), .A3(new_n642), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n910), .A2(new_n642), .A3(new_n969), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G204gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(G1353gat));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n300), .A3(new_n583), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n910), .A2(new_n583), .A3(new_n969), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  NAND3_X1  g786(.A1(new_n967), .A2(new_n301), .A3(new_n617), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n910), .A2(new_n617), .A3(new_n969), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n989), .B2(new_n301), .ZN(G1355gat));
endmodule


