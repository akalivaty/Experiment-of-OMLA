//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n212), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n211), .B(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n229), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  XNOR2_X1  g0041(.A(KEYINPUT3), .B(G33), .ZN(new_n242));
  INV_X1    g0042(.A(G1698), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G222), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G223), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n242), .A2(G1698), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n246), .B1(new_n247), .B2(new_n242), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT67), .A2(G45), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT67), .A2(G45), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n254), .A2(new_n255), .A3(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n253), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n255), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT67), .A2(G45), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n258), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n266), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n266), .B(KEYINPUT69), .C1(new_n267), .C2(new_n272), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n252), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G200), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n208), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n209), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G50), .A2(G58), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n209), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n281), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n270), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n281), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n270), .A2(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G50), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n295), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n291), .B(new_n298), .C1(G50), .C2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT9), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n277), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT10), .B1(new_n279), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n277), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G190), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n278), .A4(new_n301), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n277), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n300), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n294), .A2(new_n295), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n289), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n296), .A2(G68), .A3(new_n297), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n289), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n247), .B2(new_n283), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n281), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(KEYINPUT11), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(KEYINPUT11), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n316), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n329), .A2(new_n319), .A3(KEYINPUT74), .A4(new_n321), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n312), .A2(KEYINPUT75), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n272), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n271), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G238), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n266), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n242), .A2(G232), .A3(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(new_n341), .C1(new_n244), .C2(new_n267), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n251), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n334), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  AND4_X1   g0144(.A1(new_n334), .A2(new_n343), .A3(new_n266), .A4(new_n338), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n332), .B(new_n333), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n266), .A3(new_n338), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT73), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT13), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n339), .B(new_n343), .C1(KEYINPUT73), .C2(new_n334), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(G179), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n339), .A2(new_n334), .A3(new_n343), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n332), .B1(new_n355), .B2(new_n333), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n331), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n328), .A2(new_n330), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n349), .A2(new_n350), .A3(G190), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(G200), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G244), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n272), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n260), .B2(new_n265), .ZN(new_n364));
  INV_X1    g0164(.A(G238), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n249), .A2(new_n365), .B1(new_n203), .B2(new_n242), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n245), .A2(KEYINPUT71), .A3(G232), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT71), .ZN(new_n368));
  INV_X1    g0168(.A(G232), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n244), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n364), .B1(new_n371), .B2(new_n269), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n312), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n310), .B(new_n364), .C1(new_n371), .C2(new_n269), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n296), .A2(G77), .A3(new_n297), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G20), .A2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n283), .ZN(new_n378));
  INV_X1    g0178(.A(new_n282), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n285), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n281), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n375), .B1(G77), .B2(new_n299), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n374), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n372), .B2(G200), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n302), .B2(new_n372), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n357), .A2(new_n361), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT80), .ZN(new_n387));
  AND2_X1   g0187(.A1(KEYINPUT3), .A2(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT3), .A2(G33), .ZN(new_n389));
  OAI211_X1 g0189(.A(G226), .B(G1698), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n248), .A2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT77), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(G33), .A3(G87), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(new_n392), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT78), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n242), .A2(new_n391), .B1(new_n394), .B2(new_n396), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(new_n390), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n269), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n269), .A2(G232), .A3(new_n271), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n266), .A2(new_n302), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n387), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n266), .A2(new_n405), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n401), .B1(new_n400), .B2(new_n390), .ZN(new_n411));
  AND4_X1   g0211(.A1(new_n401), .A2(new_n390), .A3(new_n392), .A4(new_n397), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n251), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(G190), .B(new_n404), .C1(new_n260), .C2(new_n265), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT80), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n407), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n282), .B1(new_n270), .B2(G20), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n296), .A2(new_n417), .B1(new_n317), .B2(new_n282), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT3), .ZN(new_n421));
  INV_X1    g0221(.A(G33), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(KEYINPUT3), .A2(G33), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n209), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n423), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n424), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n289), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G58), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n289), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G58), .A2(G68), .ZN(new_n432));
  OAI21_X1  g0232(.A(G20), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G159), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n286), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n420), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(new_n281), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n388), .A2(new_n389), .A3(new_n426), .A4(G20), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n289), .B1(new_n438), .B2(KEYINPUT76), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT76), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n427), .A2(new_n440), .A3(new_n428), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n419), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n416), .A2(new_n444), .A3(KEYINPUT17), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT17), .B1(new_n416), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G169), .B1(new_n403), .B2(new_n409), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n404), .B1(new_n260), .B2(new_n265), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n413), .A2(G179), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n436), .A2(new_n281), .ZN(new_n452));
  AOI211_X1 g0252(.A(new_n420), .B(new_n435), .C1(new_n439), .C2(new_n441), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n418), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT79), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n451), .A2(new_n454), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT18), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT79), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n447), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n315), .A2(new_n386), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(KEYINPUT89), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n242), .A2(new_n209), .A3(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(KEYINPUT89), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n242), .A2(new_n471), .A3(new_n209), .A4(G87), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n209), .B2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n475), .A2(new_n476), .B1(new_n478), .B2(new_n209), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(KEYINPUT24), .A3(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n281), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT90), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n294), .A2(new_n203), .A3(new_n295), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT25), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n317), .A2(KEYINPUT90), .A3(KEYINPUT25), .A4(new_n203), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT91), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n486), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n486), .B2(new_n487), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n488), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n270), .A2(G33), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n296), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT92), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n493), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n484), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT5), .B(G41), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G1), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G264), .A3(new_n269), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(new_n269), .A3(G274), .A4(new_n503), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G257), .B(G1698), .C1(new_n388), .C2(new_n389), .ZN(new_n508));
  OAI211_X1 g0308(.A(G250), .B(new_n243), .C1(new_n388), .C2(new_n389), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT93), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n269), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT93), .A4(new_n510), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n310), .B2(new_n515), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n500), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT20), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n209), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n202), .A2(KEYINPUT81), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT81), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n525), .B2(new_n422), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n280), .A2(new_n208), .B1(G20), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n519), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT81), .B(G97), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G33), .ZN(new_n532));
  OAI211_X1 g0332(.A(KEYINPUT20), .B(new_n528), .C1(new_n532), .C2(new_n521), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n296), .A2(KEYINPUT88), .A3(G116), .A4(new_n494), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n299), .A2(G116), .A3(new_n381), .A4(new_n494), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT88), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n317), .A2(new_n527), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(G1698), .C1(new_n388), .C2(new_n389), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(new_n243), .C1(new_n388), .C2(new_n389), .ZN(new_n542));
  XOR2_X1   g0342(.A(KEYINPUT87), .B(G303), .Z(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n242), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n251), .B1(new_n503), .B2(new_n501), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n544), .A2(new_n251), .B1(new_n545), .B2(G270), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n312), .B1(new_n546), .B2(new_n506), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n506), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(new_n310), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n549), .A2(new_n551), .B1(new_n540), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n302), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n408), .B1(new_n546), .B2(new_n506), .ZN(new_n556));
  OR3_X1    g0356(.A1(new_n555), .A2(new_n540), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n513), .A2(new_n514), .ZN(new_n558));
  INV_X1    g0358(.A(new_n507), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n302), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n515), .B2(G200), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n484), .C1(new_n498), .C2(new_n499), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n518), .A2(new_n554), .A3(new_n557), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n504), .A2(G257), .A3(new_n269), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n506), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(KEYINPUT4), .A2(G244), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n243), .B(new_n567), .C1(new_n388), .C2(new_n389), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n362), .B1(new_n423), .B2(new_n424), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n520), .C1(new_n569), .C2(KEYINPUT4), .ZN(new_n570));
  OAI21_X1  g0370(.A(G250), .B1(new_n388), .B2(new_n389), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n243), .B1(new_n571), .B2(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n251), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n573), .A3(new_n302), .ZN(new_n574));
  OAI21_X1  g0374(.A(G244), .B1(new_n388), .B2(new_n389), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(G33), .B2(G283), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n242), .B2(G250), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n568), .C1(new_n243), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n565), .B1(new_n579), .B2(new_n251), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n574), .B1(new_n580), .B2(G200), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n317), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(new_n495), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(G97), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n427), .A2(new_n428), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G107), .B1(G77), .B2(new_n285), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT82), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G97), .A2(G107), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n204), .A2(KEYINPUT82), .A3(new_n590), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n203), .A2(KEYINPUT6), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n522), .B2(new_n524), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G20), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n586), .B(new_n381), .C1(new_n588), .C2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n388), .A2(new_n389), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT7), .B1(new_n603), .B2(new_n209), .ZN(new_n604));
  OAI21_X1  g0404(.A(G107), .B1(new_n604), .B2(new_n438), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n285), .A2(G77), .ZN(new_n606));
  XNOR2_X1  g0406(.A(G97), .B(G107), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT6), .B1(new_n607), .B2(new_n589), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n598), .B1(new_n608), .B2(new_n594), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n605), .B(new_n606), .C1(new_n609), .C2(new_n209), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT83), .B1(new_n610), .B2(new_n281), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n581), .B(new_n585), .C1(new_n602), .C2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n531), .B2(new_n283), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G87), .A2(G107), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n522), .A2(new_n524), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n209), .B1(new_n341), .B2(new_n613), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n242), .A2(new_n209), .A3(G68), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n281), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n317), .A2(new_n377), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n296), .A2(G87), .A3(new_n494), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n365), .A2(new_n243), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n362), .A2(G1698), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n625), .B(new_n626), .C1(new_n388), .C2(new_n389), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n269), .B1(new_n627), .B2(new_n477), .ZN(new_n628));
  INV_X1    g0428(.A(G250), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n257), .B1(new_n629), .B2(KEYINPUT84), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n503), .ZN(new_n631));
  OAI211_X1 g0431(.A(KEYINPUT84), .B(G250), .C1(new_n502), .C2(G1), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n251), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  AOI21_X1  g0435(.A(G274), .B1(new_n635), .B2(G250), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n270), .A2(G45), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n269), .ZN(new_n639));
  NOR2_X1   g0439(.A1(G238), .A2(G1698), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n362), .B2(G1698), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n478), .B1(new_n641), .B2(new_n242), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n639), .B(G190), .C1(new_n642), .C2(new_n269), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n624), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(G169), .B1(new_n628), .B2(new_n633), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n639), .B(G179), .C1(new_n642), .C2(new_n269), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n620), .A2(new_n281), .B1(new_n317), .B2(new_n377), .ZN(new_n650));
  INV_X1    g0450(.A(new_n377), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n495), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT85), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n645), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n610), .A2(new_n281), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n586), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n610), .A2(KEYINPUT83), .A3(new_n281), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n584), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n580), .A2(new_n310), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n566), .A2(new_n573), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n312), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n612), .B(new_n655), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT86), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n585), .B1(new_n602), .B2(new_n611), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n660), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT86), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n612), .A4(new_n655), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n563), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n465), .A2(new_n671), .ZN(G372));
  INV_X1    g0472(.A(new_n314), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT94), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n383), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n373), .A2(KEYINPUT94), .A3(new_n374), .A4(new_n382), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n357), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n447), .A2(new_n361), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n460), .B(new_n462), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n673), .B1(new_n680), .B2(new_n309), .ZN(new_n681));
  INV_X1    g0481(.A(new_n465), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n650), .A2(new_n652), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n648), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n655), .A2(new_n666), .A3(new_n667), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n659), .A2(new_n663), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n685), .A2(new_n645), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n553), .A2(new_n540), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n540), .A2(new_n547), .A3(new_n550), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n550), .B1(new_n540), .B2(new_n547), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n500), .B2(new_n517), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n668), .A2(new_n562), .A3(new_n612), .A4(new_n690), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n687), .B(new_n691), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n681), .B1(new_n682), .B2(new_n699), .ZN(G369));
  NAND3_X1  g0500(.A1(new_n270), .A2(new_n209), .A3(G13), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G343), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT95), .Z(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n540), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n554), .A2(new_n557), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n695), .A2(new_n540), .A3(new_n706), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n706), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n500), .A2(new_n517), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n500), .A2(new_n706), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n562), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n716), .B1(new_n518), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n554), .A2(new_n706), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n716), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n213), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G41), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G1), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n531), .A2(new_n527), .A3(new_n615), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n727), .A2(new_n728), .B1(new_n206), .B2(new_n726), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n688), .A2(new_n689), .A3(new_n655), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n690), .A2(new_n666), .A3(new_n667), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n684), .C1(new_n689), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n696), .A2(new_n697), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT29), .B(new_n714), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n699), .A2(new_n706), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n665), .A2(new_n670), .ZN(new_n738));
  INV_X1    g0538(.A(new_n563), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n714), .ZN(new_n740));
  INV_X1    g0540(.A(new_n647), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n580), .A2(new_n515), .A3(new_n741), .A4(new_n546), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n741), .A2(new_n546), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(KEYINPUT30), .A3(new_n580), .A4(new_n515), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n639), .B1(new_n642), .B2(new_n269), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n552), .A2(new_n661), .A3(new_n310), .A4(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n744), .B(new_n746), .C1(new_n748), .C2(new_n515), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n706), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n737), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n730), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(new_n712), .A2(G330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n209), .A2(G13), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n270), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OR3_X1    g0565(.A1(new_n765), .A2(new_n725), .A3(KEYINPUT97), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT97), .B1(new_n765), .B2(new_n725), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n713), .A2(new_n761), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT98), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n208), .B1(G20), .B2(new_n312), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n209), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G87), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n773), .A2(new_n302), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n209), .A2(new_n310), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n776), .B1(new_n203), .B2(new_n777), .C1(new_n781), .C2(new_n289), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n773), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G159), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n778), .A2(new_n783), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n778), .A2(G190), .A3(new_n408), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n242), .B1(new_n788), .B2(new_n247), .C1(new_n430), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n779), .A2(new_n302), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G50), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n302), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n209), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n202), .B2(new_n795), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n782), .A2(new_n787), .A3(new_n790), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n795), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G294), .A2(new_n798), .B1(new_n780), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n777), .ZN(new_n802));
  INV_X1    g0602(.A(new_n789), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G322), .B1(new_n785), .B2(G329), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n603), .C1(new_n805), .C2(new_n788), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n791), .A2(G326), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n774), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n802), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n772), .B1(new_n797), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n724), .A2(new_n603), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n812), .A2(G355), .B1(new_n527), .B2(new_n724), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n237), .A2(new_n502), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n724), .A2(new_n242), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n261), .A2(new_n263), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n206), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n813), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n772), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n768), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n821), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n811), .B(new_n823), .C1(new_n712), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n771), .A2(new_n825), .ZN(G396));
  AND3_X1   g0626(.A1(new_n385), .A2(new_n383), .A3(new_n714), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n698), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT99), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT99), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n698), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n675), .A2(new_n382), .A3(new_n676), .A4(new_n706), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n706), .A2(new_n382), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n385), .A2(new_n383), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n736), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n769), .B1(new_n837), .B2(new_n757), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n757), .B2(new_n837), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n772), .A2(new_n819), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n769), .B1(G77), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n788), .A2(new_n527), .B1(new_n784), .B2(new_n805), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n242), .B(new_n842), .C1(G294), .C2(new_n803), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n775), .A2(G107), .ZN(new_n844));
  INV_X1    g0644(.A(new_n777), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n791), .A2(G303), .B1(new_n845), .B2(G87), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G97), .A2(new_n798), .B1(new_n780), .B2(G283), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n843), .A2(new_n844), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n788), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n803), .A2(G143), .B1(new_n849), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n781), .B2(new_n284), .C1(new_n851), .C2(new_n792), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT34), .Z(new_n853));
  AOI22_X1  g0653(.A1(new_n798), .A2(G58), .B1(new_n775), .B2(G50), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n845), .A2(G68), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n603), .B1(new_n785), .B2(G132), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n848), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n841), .B1(new_n858), .B2(new_n772), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n820), .B2(new_n836), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n839), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  OR2_X1    g0662(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(G116), .A3(new_n210), .A4(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT36), .Z(new_n866));
  OAI211_X1 g0666(.A(new_n207), .B(G77), .C1(new_n430), .C2(new_n289), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n793), .A2(G68), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n270), .B(G13), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n331), .A2(new_n706), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n357), .A2(new_n361), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n357), .B2(new_n361), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n383), .A2(new_n706), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT100), .Z(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n832), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n443), .A2(new_n281), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n418), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n704), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n464), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n451), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n416), .A2(new_n444), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n454), .B1(new_n451), .B2(new_n704), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n884), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n464), .A2(new_n882), .B1(new_n891), .B2(new_n888), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n460), .A2(new_n462), .ZN(new_n896));
  INV_X1    g0696(.A(new_n704), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n877), .A2(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n889), .A2(new_n886), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT101), .B1(new_n901), .B2(new_n890), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n890), .B1(new_n889), .B2(new_n886), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT101), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n905), .A3(new_n891), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n444), .A2(new_n897), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT17), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n886), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n416), .A2(new_n444), .A3(KEYINPUT17), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(new_n896), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT102), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n905), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n891), .B1(new_n903), .B2(new_n904), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n884), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT102), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(new_n899), .A4(new_n893), .ZN(new_n920));
  INV_X1    g0720(.A(new_n893), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n888), .A2(new_n891), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n883), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT39), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n914), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n357), .A2(new_n706), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n898), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n465), .B(new_n735), .C1(new_n736), .C2(KEYINPUT29), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n681), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n833), .A2(new_n835), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n357), .A2(new_n361), .ZN(new_n934));
  INV_X1    g0734(.A(new_n871), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n357), .A2(new_n361), .A3(new_n871), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n895), .A2(new_n756), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n754), .B1(new_n671), .B2(new_n714), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n836), .B1(new_n872), .B2(new_n873), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n941), .A2(new_n942), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n918), .A2(new_n893), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n939), .A2(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n682), .B2(new_n941), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n465), .A3(new_n756), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n270), .B2(new_n763), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n932), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n870), .B1(new_n951), .B2(new_n952), .ZN(G367));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n668), .B(new_n612), .C1(new_n659), .C2(new_n714), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n688), .A2(new_n706), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n722), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT45), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n722), .A2(new_n957), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT44), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n959), .A2(new_n720), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n720), .B1(new_n959), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n719), .B(new_n721), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n712), .A2(KEYINPUT104), .A3(G330), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n966), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n758), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n725), .B(KEYINPUT41), .Z(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT105), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n970), .A2(new_n758), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n959), .A2(new_n720), .A3(new_n961), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n959), .A2(new_n961), .ZN(new_n977));
  INV_X1    g0777(.A(new_n720), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n759), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT105), .ZN(new_n982));
  INV_X1    g0782(.A(new_n973), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n765), .B1(new_n974), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n719), .A2(new_n721), .A3(new_n957), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n668), .B1(new_n955), .B2(new_n518), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n986), .A2(KEYINPUT42), .B1(new_n714), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(KEYINPUT42), .B2(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n706), .A2(new_n624), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n690), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n684), .B2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT103), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n978), .A2(new_n957), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n996), .B2(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n996), .A2(new_n998), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n954), .B1(new_n985), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(new_n1005));
  AOI211_X1 g0805(.A(KEYINPUT105), .B(new_n973), .C1(new_n980), .C2(new_n759), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n764), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1003), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(KEYINPUT106), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n795), .A2(new_n289), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G58), .B2(new_n775), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n434), .B2(new_n781), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n803), .A2(G150), .B1(new_n785), .B2(G137), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n242), .C1(new_n793), .C2(new_n788), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n845), .A2(G77), .ZN(new_n1016));
  INV_X1    g0816(.A(G143), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n792), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1013), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT110), .Z(new_n1020));
  NAND3_X1  g0820(.A1(new_n775), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT108), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G107), .A2(new_n798), .B1(new_n780), .B2(G294), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT109), .B(G317), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n788), .A2(new_n801), .B1(new_n784), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n543), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n242), .B(new_n1025), .C1(new_n1026), .C2(new_n803), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n791), .A2(G311), .B1(new_n845), .B2(new_n525), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n774), .B2(new_n527), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1023), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1022), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n772), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n233), .A2(new_n815), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n822), .C1(new_n213), .C2(new_n377), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT107), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n768), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1034), .B(new_n1040), .C1(new_n824), .C2(new_n992), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1010), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT111), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n971), .A2(new_n765), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n242), .B1(new_n785), .B2(G326), .ZN(new_n1045));
  INV_X1    g0845(.A(G294), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n795), .A2(new_n801), .B1(new_n774), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1024), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n803), .A2(new_n1048), .B1(new_n1026), .B2(new_n849), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n791), .A2(G322), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n805), .C2(new_n781), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1045), .B1(new_n527), .B2(new_n777), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n603), .B1(new_n785), .B2(G150), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n247), .B2(new_n774), .C1(new_n202), .C2(new_n777), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT112), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n798), .A2(new_n651), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n793), .B2(new_n789), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT113), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n781), .A2(new_n282), .B1(new_n788), .B2(new_n289), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G159), .B2(new_n791), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT114), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n772), .B1(new_n1057), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n815), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n229), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n816), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n728), .B2(new_n812), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n379), .A2(new_n793), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n502), .B1(new_n289), .B2(new_n247), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1074), .A2(new_n728), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1072), .A2(new_n1076), .B1(G107), .B2(new_n213), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n768), .B1(new_n1077), .B2(new_n822), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1068), .B(new_n1078), .C1(new_n719), .C2(new_n824), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1044), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n975), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n970), .A2(new_n758), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n725), .B(KEYINPUT115), .Z(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1080), .A2(new_n1084), .ZN(G393));
  NAND3_X1  g0885(.A1(new_n955), .A2(new_n956), .A3(new_n821), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n822), .B1(new_n213), .B2(new_n531), .C1(new_n240), .C2(new_n1069), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n769), .A2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n792), .A2(new_n284), .B1(new_n434), .B2(new_n789), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  NOR2_X1   g0890(.A1(new_n795), .A2(new_n247), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G68), .B2(new_n775), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n242), .B1(new_n784), .B2(new_n1017), .C1(new_n282), .C2(new_n788), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n780), .A2(G50), .B1(new_n845), .B2(G87), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G317), .A2(new_n791), .B1(new_n803), .B2(G311), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n603), .B1(new_n788), .B2(new_n1046), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G322), .B2(new_n785), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n798), .A2(G116), .B1(new_n845), .B2(G107), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n780), .A2(new_n1026), .B1(new_n775), .B2(G283), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1090), .A2(new_n1096), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1088), .B1(new_n1104), .B2(new_n772), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n964), .A2(new_n765), .B1(new_n1086), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n980), .A2(new_n1083), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n964), .A2(new_n975), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(G390));
  OAI21_X1  g0909(.A(new_n714), .B1(new_n733), .B2(new_n734), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n876), .B1(new_n1110), .B2(new_n933), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n874), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n926), .A3(new_n944), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n698), .A2(new_n830), .A3(new_n827), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n830), .B1(new_n698), .B2(new_n827), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n876), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n927), .B1(new_n1117), .B2(new_n1112), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1114), .B1(new_n925), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G330), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n941), .A2(new_n874), .A3(new_n1120), .A4(new_n933), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n740), .B2(new_n755), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n836), .A3(new_n1112), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n1114), .C1(new_n925), .C2(new_n1118), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n765), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n769), .B1(new_n379), .B2(new_n840), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n788), .A2(new_n1128), .B1(new_n784), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n603), .B(new_n1130), .C1(G132), .C2(new_n803), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n774), .A2(new_n284), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n791), .A2(G128), .B1(new_n845), .B2(G50), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G159), .A2(new_n798), .B1(new_n780), .B2(G137), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n788), .A2(new_n531), .B1(new_n784), .B2(new_n1046), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n242), .B(new_n1137), .C1(G116), .C2(new_n803), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n776), .A3(new_n855), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1091), .B1(G283), .B2(new_n791), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n203), .B2(new_n781), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1127), .B1(new_n1142), .B2(new_n772), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n925), .B2(new_n820), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1126), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT117), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1126), .A2(KEYINPUT117), .A3(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n930), .B(new_n681), .C1(new_n682), .C2(new_n757), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1112), .B1(new_n1123), .B2(new_n836), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1111), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1124), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1117), .B1(new_n1121), .B2(new_n1151), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n918), .A2(new_n899), .A3(new_n893), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(KEYINPUT102), .B1(new_n895), .B2(KEYINPUT39), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n920), .C1(new_n877), .C2(new_n927), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1124), .B1(new_n1160), .B2(new_n1114), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1125), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1122), .A2(new_n1125), .A3(new_n1156), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1083), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT116), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(KEYINPUT116), .A3(new_n1083), .A4(new_n1164), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1149), .A2(new_n1167), .A3(new_n1168), .ZN(G378));
  AOI21_X1  g0969(.A(new_n673), .B1(new_n308), .B2(new_n304), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n300), .A2(new_n704), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n315), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1172), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n945), .B2(G330), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n883), .A2(new_n922), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1182), .A2(new_n884), .B1(new_n883), .B2(new_n892), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n756), .A2(new_n938), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n940), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n943), .A2(new_n944), .ZN(new_n1186));
  AND4_X1   g0986(.A1(G330), .A2(new_n1185), .A3(new_n1186), .A4(new_n1180), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n929), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(G330), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1180), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1185), .A2(new_n1186), .A3(G330), .A4(new_n1180), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1191), .A2(new_n928), .A3(new_n898), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1188), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n765), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n769), .B1(G50), .B2(new_n840), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT119), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n202), .A2(new_n781), .B1(new_n792), .B2(new_n527), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1011), .B(new_n1198), .C1(G77), .C2(new_n775), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n603), .A2(new_n262), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n651), .B2(new_n849), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(new_n801), .C2(new_n784), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n803), .A2(KEYINPUT118), .A3(G107), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT118), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n789), .B2(new_n203), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n430), .C2(new_n777), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT58), .ZN(new_n1208));
  INV_X1    g1008(.A(G132), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1129), .A2(new_n792), .B1(new_n781), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n803), .A2(G128), .B1(new_n849), .B2(G137), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n774), .B2(new_n1128), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G150), .C2(new_n798), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n845), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1207), .A2(KEYINPUT58), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1200), .B(new_n793), .C1(G33), .C2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1208), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1197), .B1(new_n1222), .B2(new_n772), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1180), .B2(new_n820), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1195), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1150), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1164), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1194), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1083), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n1227), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1225), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G375));
  NAND2_X1  g1035(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n1226), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT120), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1238), .A2(new_n973), .A3(new_n1156), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n765), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n769), .B1(G68), .B2(new_n840), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n792), .A2(new_n1209), .B1(new_n774), .B2(new_n434), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G50), .B2(new_n798), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n603), .B1(new_n785), .B2(G128), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n803), .A2(G137), .B1(new_n849), .B2(G150), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1128), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n780), .A2(new_n1246), .B1(new_n845), .B2(G58), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n603), .B1(new_n789), .B2(new_n801), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G303), .B2(new_n785), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n791), .A2(G294), .B1(new_n775), .B2(G97), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1016), .A3(new_n1061), .A4(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n780), .A2(G116), .B1(new_n849), .B2(G107), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT121), .Z(new_n1254));
  OAI21_X1  g1054(.A(new_n1248), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1255), .B2(new_n772), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1112), .B2(new_n820), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1257), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT122), .Z(new_n1259));
  NAND2_X1  g1059(.A1(new_n1239), .A2(new_n1259), .ZN(G381));
  XOR2_X1   g1060(.A(new_n1234), .B(KEYINPUT123), .Z(new_n1261));
  AND3_X1   g1061(.A1(new_n1165), .A2(new_n1126), .A3(new_n1144), .ZN(new_n1262));
  INV_X1    g1062(.A(G396), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1080), .A2(new_n1084), .A3(new_n1263), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(G381), .A2(G384), .A3(G390), .A4(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1261), .A2(new_n1262), .A3(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(G387), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT124), .ZN(G407));
  INV_X1    g1068(.A(G213), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(G343), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1262), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1261), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G407), .A2(new_n1272), .ZN(G409));
  OAI211_X1 g1073(.A(new_n1195), .B(new_n1224), .C1(new_n1228), .C2(new_n973), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1262), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1234), .A2(KEYINPUT125), .A3(G378), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT125), .B1(new_n1234), .B2(G378), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1270), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1231), .B1(new_n1237), .B2(KEYINPUT60), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1157), .A2(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1238), .B2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1282), .A2(new_n1259), .A3(G384), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1282), .B2(new_n1259), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n1279), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G2897), .B(new_n1270), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1282), .A2(new_n1259), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n861), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1282), .A2(new_n1259), .A3(G384), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(G2897), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1234), .A2(G378), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1234), .A2(G378), .A3(KEYINPUT125), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1298), .A2(new_n1299), .B1(new_n1262), .B2(new_n1274), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1295), .B1(new_n1300), .B2(new_n1270), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1278), .A2(new_n1302), .A3(new_n1279), .A4(new_n1285), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1287), .A2(new_n1288), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1264), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1263), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1306));
  OAI21_X1  g1106(.A(G390), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT111), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1306), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1264), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1307), .B1(new_n1310), .B2(G390), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1010), .A2(new_n1041), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1010), .B2(new_n1041), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1311), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1042), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT126), .B1(new_n1318), .B2(new_n1312), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1304), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1295), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1286), .A2(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1279), .A4(new_n1285), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1321), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT127), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1321), .A2(KEYINPUT127), .A3(new_n1328), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(G405));
  NAND2_X1  g1133(.A1(G375), .A2(new_n1262), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1335), .B(new_n1285), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1320), .B(new_n1336), .ZN(G402));
endmodule


