

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XNOR2_X1 U325 ( .A(n451), .B(n450), .ZN(n532) );
  XOR2_X1 U326 ( .A(n322), .B(n352), .Z(n293) );
  XNOR2_X1 U327 ( .A(KEYINPUT25), .B(KEYINPUT94), .ZN(n467) );
  XNOR2_X1 U328 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U329 ( .A(KEYINPUT111), .ZN(n396) );
  INV_X1 U330 ( .A(KEYINPUT54), .ZN(n417) );
  INV_X1 U331 ( .A(G127GAT), .ZN(n296) );
  XNOR2_X1 U332 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U333 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n475) );
  XNOR2_X1 U334 ( .A(n299), .B(n298), .ZN(n447) );
  XNOR2_X1 U335 ( .A(n476), .B(n475), .ZN(n516) );
  INV_X1 U336 ( .A(G190GAT), .ZN(n454) );
  XNOR2_X1 U337 ( .A(n453), .B(KEYINPUT118), .ZN(n568) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n479) );
  XNOR2_X1 U339 ( .A(KEYINPUT92), .B(n470), .ZN(n546) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U341 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U342 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT77), .B(KEYINPUT0), .Z(n295) );
  XNOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT76), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n299) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G120GAT), .ZN(n297) );
  XOR2_X1 U348 ( .A(KEYINPUT87), .B(KEYINPUT89), .Z(n301) );
  XNOR2_X1 U349 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U351 ( .A(KEYINPUT88), .B(n302), .Z(n304) );
  NAND2_X1 U352 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U354 ( .A(n305), .B(KEYINPUT1), .Z(n311) );
  XOR2_X1 U355 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n307) );
  XNOR2_X1 U356 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(n308), .ZN(n436) );
  INV_X1 U359 ( .A(n436), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n309), .B(KEYINPUT90), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U362 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n313) );
  XOR2_X1 U363 ( .A(G29GAT), .B(G85GAT), .Z(n322) );
  XOR2_X1 U364 ( .A(G148GAT), .B(G57GAT), .Z(n359) );
  XNOR2_X1 U365 ( .A(n322), .B(n359), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n315), .B(n314), .Z(n317) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G162GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n447), .B(n318), .ZN(n470) );
  INV_X1 U371 ( .A(KEYINPUT47), .ZN(n392) );
  XOR2_X1 U372 ( .A(G36GAT), .B(G218GAT), .Z(n403) );
  XOR2_X1 U373 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  XOR2_X1 U374 ( .A(n403), .B(n424), .Z(n320) );
  XNOR2_X1 U375 ( .A(G99GAT), .B(G106GAT), .ZN(n319) );
  XOR2_X1 U376 ( .A(n320), .B(n319), .Z(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n321), .B(KEYINPUT70), .ZN(n352) );
  NAND2_X1 U379 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n293), .B(n323), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n327) );
  XNOR2_X1 U382 ( .A(G190GAT), .B(G134GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n335) );
  XOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n329) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G92GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n331) );
  XNOR2_X1 U388 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n542) );
  INV_X1 U392 ( .A(n542), .ZN(n558) );
  XOR2_X1 U393 ( .A(KEYINPUT69), .B(G113GAT), .Z(n337) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(G197GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n356) );
  XOR2_X1 U396 ( .A(G43GAT), .B(G15GAT), .Z(n444) );
  INV_X1 U397 ( .A(G50GAT), .ZN(n338) );
  NAND2_X1 U398 ( .A1(G141GAT), .A2(n338), .ZN(n341) );
  INV_X1 U399 ( .A(G141GAT), .ZN(n339) );
  NAND2_X1 U400 ( .A1(n339), .A2(G50GAT), .ZN(n340) );
  NAND2_X1 U401 ( .A1(n341), .A2(n340), .ZN(n343) );
  XNOR2_X1 U402 ( .A(G29GAT), .B(G36GAT), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U404 ( .A(n444), .B(n344), .Z(n346) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n348) );
  XNOR2_X1 U408 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U410 ( .A(n350), .B(n349), .Z(n354) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G1GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n351), .B(G8GAT), .ZN(n375) );
  XNOR2_X1 U413 ( .A(n352), .B(n375), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U415 ( .A(n356), .B(n355), .Z(n548) );
  XOR2_X1 U416 ( .A(KEYINPUT72), .B(G85GAT), .Z(n358) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(G120GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n363) );
  XOR2_X1 U420 ( .A(G99GAT), .B(G71GAT), .Z(n440) );
  XNOR2_X1 U421 ( .A(G106GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n361), .B(G204GAT), .ZN(n431) );
  XNOR2_X1 U423 ( .A(n440), .B(n431), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n370) );
  XOR2_X1 U425 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n365) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U428 ( .A(n366), .B(KEYINPUT31), .Z(n368) );
  XOR2_X1 U429 ( .A(G92GAT), .B(G64GAT), .Z(n406) );
  XOR2_X1 U430 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n374) );
  XNOR2_X1 U431 ( .A(n406), .B(n374), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n580) );
  XNOR2_X1 U434 ( .A(KEYINPUT41), .B(n580), .ZN(n551) );
  NAND2_X1 U435 ( .A1(n548), .A2(n551), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n371), .B(KEYINPUT46), .ZN(n389) );
  XOR2_X1 U437 ( .A(G211GAT), .B(G71GAT), .Z(n373) );
  XNOR2_X1 U438 ( .A(G15GAT), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n388) );
  XOR2_X1 U440 ( .A(n374), .B(G78GAT), .Z(n377) );
  XNOR2_X1 U441 ( .A(n375), .B(G155GAT), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n379) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U446 ( .A(n381), .B(n380), .Z(n386) );
  XOR2_X1 U447 ( .A(KEYINPUT75), .B(G64GAT), .Z(n383) );
  XNOR2_X1 U448 ( .A(G127GAT), .B(G57GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n384), .B(KEYINPUT15), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n583) );
  NAND2_X1 U453 ( .A1(n389), .A2(n583), .ZN(n390) );
  NOR2_X1 U454 ( .A1(n558), .A2(n390), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n399) );
  XNOR2_X1 U456 ( .A(KEYINPUT36), .B(n542), .ZN(n589) );
  NOR2_X1 U457 ( .A1(n589), .A2(n583), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n393), .B(KEYINPUT45), .ZN(n394) );
  NAND2_X1 U459 ( .A1(n394), .A2(n580), .ZN(n395) );
  NOR2_X1 U460 ( .A1(n395), .A2(n548), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  NOR2_X1 U462 ( .A1(n399), .A2(n398), .ZN(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT48), .B(n400), .ZN(n530) );
  XOR2_X1 U464 ( .A(G211GAT), .B(KEYINPUT21), .Z(n402) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(KEYINPUT84), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n430) );
  XOR2_X1 U467 ( .A(n403), .B(n430), .Z(n405) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U470 ( .A(n407), .B(n406), .Z(n409) );
  XNOR2_X1 U471 ( .A(G8GAT), .B(G204GAT), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n416) );
  XOR2_X1 U473 ( .A(G176GAT), .B(G183GAT), .Z(n411) );
  XNOR2_X1 U474 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U476 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n413) );
  XNOR2_X1 U477 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U479 ( .A(n415), .B(n414), .Z(n451) );
  XNOR2_X1 U480 ( .A(n416), .B(n451), .ZN(n518) );
  INV_X1 U481 ( .A(n518), .ZN(n459) );
  NOR2_X1 U482 ( .A1(n530), .A2(n459), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n419), .B(KEYINPUT116), .ZN(n420) );
  NOR2_X1 U485 ( .A1(n546), .A2(n420), .ZN(n573) );
  XOR2_X1 U486 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n422) );
  XNOR2_X1 U487 ( .A(G218GAT), .B(KEYINPUT23), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U489 ( .A(n423), .B(G148GAT), .Z(n426) );
  XNOR2_X1 U490 ( .A(G22GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT83), .B(KEYINPUT24), .Z(n428) );
  NAND2_X1 U493 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U495 ( .A(n429), .B(KEYINPUT22), .Z(n433) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n465) );
  NAND2_X1 U500 ( .A1(n573), .A2(n465), .ZN(n439) );
  XOR2_X1 U501 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT78), .B(n440), .Z(n442) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U506 ( .A(n443), .B(KEYINPUT79), .Z(n449) );
  XNOR2_X1 U507 ( .A(n444), .B(KEYINPUT64), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n445), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U511 ( .A1(n452), .A2(n532), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n568), .A2(n542), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n548), .A2(n580), .ZN(n487) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n458) );
  XNOR2_X1 U516 ( .A(n465), .B(n458), .ZN(n525) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n525), .A2(n463), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n546), .A2(n460), .ZN(n531) );
  XOR2_X1 U520 ( .A(KEYINPUT81), .B(n532), .Z(n461) );
  NOR2_X1 U521 ( .A1(n531), .A2(n461), .ZN(n473) );
  NOR2_X1 U522 ( .A1(n465), .A2(n532), .ZN(n462) );
  XOR2_X1 U523 ( .A(n462), .B(KEYINPUT26), .Z(n571) );
  NOR2_X1 U524 ( .A1(n463), .A2(n571), .ZN(n545) );
  AND2_X1 U525 ( .A1(n532), .A2(n518), .ZN(n464) );
  XNOR2_X1 U526 ( .A(KEYINPUT93), .B(n464), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n466), .A2(n465), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n545), .A2(n469), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n485) );
  NOR2_X1 U531 ( .A1(n589), .A2(n485), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n583), .A2(n474), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n487), .A2(n516), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT38), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT100), .B(n478), .ZN(n502) );
  NAND2_X1 U536 ( .A1(n502), .A2(n532), .ZN(n482) );
  XOR2_X1 U537 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n480) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  NOR2_X1 U539 ( .A1(n558), .A2(n583), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  NOR2_X1 U541 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U542 ( .A(KEYINPUT95), .B(n486), .ZN(n505) );
  NOR2_X1 U543 ( .A1(n487), .A2(n505), .ZN(n495) );
  NAND2_X1 U544 ( .A1(n546), .A2(n495), .ZN(n488) );
  XNOR2_X1 U545 ( .A(n489), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n518), .A2(n495), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT35), .B(KEYINPUT97), .Z(n492) );
  NAND2_X1 U549 ( .A1(n495), .A2(n532), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT96), .Z(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n525), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U556 ( .A1(n502), .A2(n546), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT101), .Z(n501) );
  NAND2_X1 U560 ( .A1(n502), .A2(n518), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U563 ( .A1(n502), .A2(n525), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n507) );
  INV_X1 U566 ( .A(n548), .ZN(n574) );
  NAND2_X1 U567 ( .A1(n551), .A2(n574), .ZN(n515) );
  NOR2_X1 U568 ( .A1(n505), .A2(n515), .ZN(n511) );
  NAND2_X1 U569 ( .A1(n511), .A2(n546), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NAND2_X1 U572 ( .A1(n518), .A2(n511), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n532), .A2(n511), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U577 ( .A1(n511), .A2(n525), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n546), .A2(n526), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U584 ( .A1(n526), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U588 ( .A1(n526), .A2(n532), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n531), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n541) );
  NOR2_X1 U597 ( .A1(n574), .A2(n541), .ZN(n534) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  INV_X1 U599 ( .A(n551), .ZN(n565) );
  NOR2_X1 U600 ( .A1(n565), .A2(n541), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(n537), .ZN(G1341GAT) );
  NOR2_X1 U604 ( .A1(n583), .A2(n541), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n530), .A2(n547), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n559), .A2(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT114), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT115), .Z(n553) );
  NAND2_X1 U617 ( .A1(n559), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .Z(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  INV_X1 U621 ( .A(n583), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n559), .A2(n556), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n568), .A2(n574), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n568), .A2(n565), .ZN(n566) );
  XOR2_X1 U633 ( .A(n567), .B(n566), .Z(G1349GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n583), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  INV_X1 U637 ( .A(n571), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n588) );
  NOR2_X1 U639 ( .A1(n574), .A2(n588), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT123), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n588), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n588), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n587) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U655 ( .A(n591), .B(n590), .Z(G1355GAT) );
endmodule

