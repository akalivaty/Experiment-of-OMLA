//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(G128), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n198), .A3(new_n194), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n195), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n196), .A2(new_n198), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G143), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n200), .A3(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G131), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n214), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n212), .A2(G137), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT2), .A3(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(KEYINPUT2), .B2(G113), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n231), .A2(new_n232), .B1(KEYINPUT2), .B2(G113), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n237));
  OAI221_X1 g051(.A(new_n234), .B1(KEYINPUT2), .B2(G113), .C1(new_n231), .C2(new_n232), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(KEYINPUT68), .A3(new_n235), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n199), .A2(new_n206), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n202), .B2(new_n203), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n245), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n204), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  INV_X1    g064(.A(new_n206), .ZN(new_n251));
  INV_X1    g065(.A(new_n243), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT64), .B(G146), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n194), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n222), .A2(G131), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n218), .B1(new_n217), .B2(new_n220), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n219), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n256), .A2(new_n263), .A3(new_n260), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n242), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n244), .A2(new_n246), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n228), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(new_n241), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT28), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n228), .A2(new_n241), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n261), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n193), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n256), .A2(new_n263), .A3(new_n260), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n263), .B1(new_n256), .B2(new_n260), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n193), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(KEYINPUT72), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n228), .A2(new_n267), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n228), .B1(new_n276), .B2(new_n277), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(KEYINPUT30), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n278), .B(new_n280), .C1(new_n284), .C2(new_n241), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n286), .A2(KEYINPUT31), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n282), .ZN(new_n290));
  INV_X1    g104(.A(new_n228), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n262), .B2(new_n264), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n292), .B2(new_n281), .ZN(new_n293));
  INV_X1    g107(.A(new_n241), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(new_n278), .A3(new_n287), .A4(new_n280), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n275), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n270), .A2(new_n301), .A3(new_n274), .ZN(new_n302));
  INV_X1    g116(.A(new_n261), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT73), .B(new_n273), .C1(new_n303), .C2(new_n242), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT73), .B1(new_n272), .B2(new_n273), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n278), .B1(new_n292), .B2(new_n241), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n305), .B(new_n306), .C1(KEYINPUT28), .C2(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n302), .B(new_n193), .C1(new_n308), .C2(new_n301), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n295), .A2(new_n301), .A3(new_n278), .A4(new_n279), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n289), .A2(new_n296), .ZN(new_n315));
  INV_X1    g129(.A(new_n275), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n299), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n317), .B2(KEYINPUT32), .ZN(new_n318));
  NOR4_X1   g132(.A1(new_n297), .A2(KEYINPUT74), .A3(new_n187), .A4(new_n299), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n300), .B(new_n313), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G104), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G107), .ZN(new_n322));
  INV_X1    g136(.A(G107), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G104), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(G101), .C1(new_n325), .C2(new_n324), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n321), .A2(G107), .ZN(new_n328));
  AND2_X1   g142(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n329));
  NOR2_X1   g143(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT81), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G101), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n321), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n336), .A3(new_n322), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G116), .ZN(new_n343));
  OAI211_X1 g157(.A(G113), .B(new_n343), .C1(new_n235), .C2(new_n341), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n238), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n322), .A3(new_n337), .ZN(new_n346));
  AOI22_X1  g160(.A1(KEYINPUT4), .A2(new_n338), .B1(new_n346), .B2(G101), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n346), .A2(KEYINPUT4), .A3(G101), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n349), .B2(new_n241), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT88), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n345), .B(new_n352), .C1(new_n349), .C2(new_n241), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n210), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n266), .A2(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G224), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n364), .A3(new_n353), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n356), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n362), .B(KEYINPUT90), .Z(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n344), .A2(new_n238), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n339), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n352), .B(KEYINPUT8), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT89), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n373), .A2(KEYINPUT7), .B1(new_n361), .B2(G224), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n358), .A2(new_n359), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n368), .A2(new_n372), .A3(new_n376), .A4(new_n355), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n366), .A2(new_n310), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G210), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n366), .A2(new_n310), .A3(new_n379), .A4(new_n377), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G475), .ZN(new_n386));
  XNOR2_X1  g200(.A(G125), .B(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT16), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n357), .A2(KEYINPUT16), .A3(G140), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n195), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n189), .A2(G214), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT91), .A3(G143), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT91), .A2(G143), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT91), .A2(G143), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(G214), .A3(new_n189), .A4(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n393), .A2(new_n396), .A3(KEYINPUT17), .A4(new_n219), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n396), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n220), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n391), .B(new_n397), .C1(KEYINPUT17), .C2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n321), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT18), .A2(G131), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n398), .B(new_n403), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n207), .A2(new_n387), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n195), .B2(new_n387), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n387), .A2(new_n410), .A3(KEYINPUT19), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n387), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT93), .B1(new_n414), .B2(new_n253), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n388), .A2(G146), .A3(new_n389), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT77), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n418), .A3(new_n207), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n415), .A2(new_n417), .A3(new_n399), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n402), .B1(new_n420), .B2(new_n407), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n386), .B(new_n310), .C1(new_n409), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT20), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n420), .A2(new_n407), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n408), .B1(new_n424), .B2(new_n402), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n386), .A4(new_n310), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n402), .B1(new_n400), .B2(new_n407), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n310), .B1(new_n409), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n423), .A2(new_n427), .B1(new_n429), .B2(G475), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n194), .A2(G128), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT13), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT95), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G128), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n432), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT95), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(new_n194), .A3(KEYINPUT13), .A4(G128), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n433), .A2(new_n435), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G134), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT96), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n431), .A2(new_n435), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n212), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n444), .A3(G134), .ZN(new_n445));
  XNOR2_X1  g259(.A(G116), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT94), .B(G107), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n441), .A2(new_n443), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G116), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n450), .A2(G122), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n323), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n446), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n442), .B(new_n212), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT9), .B(G234), .Z(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT75), .B(G217), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n361), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n449), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n449), .B2(new_n455), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n310), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n463), .A2(new_n465), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n430), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(G234), .A2(G237), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n470), .A2(G952), .A3(new_n361), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT97), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n470), .A2(G902), .A3(G953), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n385), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n390), .B(G146), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n342), .A2(G128), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n342), .A2(KEYINPUT23), .A3(G128), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n481), .A2(new_n482), .B1(G119), .B2(new_n434), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G110), .ZN(new_n484));
  OR3_X1    g298(.A1(new_n434), .A2(KEYINPUT76), .A3(G119), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT76), .B1(new_n434), .B2(G119), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT24), .B(G110), .Z(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n478), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  OAI22_X1  g304(.A1(new_n483), .A2(G110), .B1(new_n487), .B2(new_n488), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n417), .A2(new_n405), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT22), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G137), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n490), .B2(new_n492), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n498), .A2(G902), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n500), .A2(KEYINPUT78), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n500), .B2(KEYINPUT78), .ZN(new_n503));
  INV_X1    g317(.A(new_n457), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(G234), .B2(new_n310), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n498), .A2(new_n499), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n505), .A2(G902), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G469), .ZN(new_n511));
  INV_X1    g325(.A(new_n260), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n203), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(G128), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n251), .B1(new_n253), .B2(new_n194), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT85), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n208), .A2(KEYINPUT83), .A3(new_n200), .A4(G128), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT85), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT83), .ZN(new_n524));
  OAI211_X1 g338(.A(G128), .B(new_n251), .C1(new_n253), .C2(new_n194), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(KEYINPUT1), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n340), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT10), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n346), .A2(G101), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT4), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n532), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n339), .B1(new_n205), .B2(new_n209), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n535), .A2(new_n256), .B1(new_n536), .B2(KEYINPUT10), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n512), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n537), .A3(new_n512), .ZN(new_n540));
  XNOR2_X1  g354(.A(G110), .B(G140), .ZN(new_n541));
  INV_X1    g355(.A(G227), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(G953), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n541), .B(new_n543), .Z(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n256), .B1(new_n347), .B2(new_n348), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(KEYINPUT10), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT10), .B1(new_n527), .B2(new_n340), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(new_n260), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n339), .A2(new_n205), .A3(new_n209), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n528), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT12), .B1(new_n260), .B2(KEYINPUT86), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n260), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n551), .B1(new_n527), .B2(new_n340), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n557), .B2(new_n512), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n550), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n545), .B1(new_n559), .B2(new_n544), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n511), .B1(new_n560), .B2(new_n310), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n555), .B1(new_n553), .B2(new_n260), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n557), .A2(new_n512), .A3(new_n554), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n540), .B(new_n544), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n544), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n550), .B2(new_n538), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n511), .A3(new_n310), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n564), .B2(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT87), .A3(new_n511), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n561), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n456), .A2(new_n310), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n574), .A2(G221), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT79), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n320), .A2(new_n477), .A3(new_n510), .A4(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n579), .B(new_n336), .Z(G3));
  INV_X1    g394(.A(new_n315), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n310), .B1(new_n581), .B2(new_n275), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n317), .B1(new_n582), .B2(G472), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n385), .A2(new_n476), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n510), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n586), .A2(new_n573), .A3(new_n577), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n430), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT33), .B1(new_n459), .B2(KEYINPUT98), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n462), .A2(new_n590), .ZN(new_n591));
  OR3_X1    g405(.A1(new_n460), .A2(new_n461), .A3(new_n590), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(G478), .A3(new_n310), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n463), .A2(new_n464), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT99), .Z(new_n597));
  NAND2_X1  g411(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n321), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT100), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT34), .ZN(G6));
  INV_X1    g415(.A(new_n468), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n423), .A2(new_n603), .A3(new_n427), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n429), .A2(G475), .ZN(new_n605));
  INV_X1    g419(.A(new_n422), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(KEYINPUT101), .A3(new_n426), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n588), .A2(new_n602), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n323), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT102), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT35), .Z(G9));
  NOR2_X1   g427(.A1(new_n589), .A2(new_n602), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n493), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n508), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n506), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n619), .A2(new_n573), .A3(new_n577), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n585), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT37), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G110), .ZN(G12));
  INV_X1    g437(.A(new_n385), .ZN(new_n624));
  INV_X1    g438(.A(G900), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n475), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n471), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n608), .A2(new_n468), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n320), .A2(new_n624), .A3(new_n620), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G128), .ZN(G30));
  XNOR2_X1  g444(.A(new_n627), .B(KEYINPUT39), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n578), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n618), .B1(new_n633), .B2(KEYINPUT40), .ZN(new_n634));
  INV_X1    g448(.A(new_n384), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n430), .A2(new_n468), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n634), .B(new_n636), .C1(KEYINPUT40), .C2(new_n633), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n383), .B(KEYINPUT38), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n295), .A2(new_n278), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n193), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n310), .B1(new_n307), .B2(new_n193), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n300), .B(new_n643), .C1(new_n318), .C2(new_n319), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n637), .A2(new_n638), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n194), .ZN(G45));
  INV_X1    g461(.A(new_n595), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n648), .A2(new_n430), .A3(new_n627), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n320), .A2(new_n624), .A3(new_n620), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  NOR2_X1   g465(.A1(new_n571), .A2(new_n511), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n575), .ZN(new_n654));
  AND4_X1   g468(.A1(KEYINPUT87), .A2(new_n567), .A3(new_n511), .A4(new_n310), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT87), .B1(new_n571), .B2(new_n511), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n653), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n320), .A2(new_n510), .A3(new_n584), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n597), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n320), .A2(new_n510), .A3(new_n584), .A4(new_n658), .ZN(new_n662));
  INV_X1    g476(.A(new_n597), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT41), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G113), .ZN(G15));
  NAND2_X1  g481(.A1(new_n609), .A2(new_n602), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n450), .ZN(G18));
  NOR3_X1   g484(.A1(new_n657), .A2(new_n619), .A3(new_n385), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n469), .A2(new_n476), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n320), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G119), .ZN(G21));
  NOR3_X1   g488(.A1(new_n657), .A2(new_n468), .A3(new_n430), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n308), .A2(new_n193), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n298), .B1(new_n581), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n297), .B2(G902), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n506), .A2(KEYINPUT104), .A3(new_n509), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT104), .B1(new_n506), .B2(new_n509), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n675), .A2(new_n679), .A3(new_n584), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT105), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  AND3_X1   g499(.A1(new_n677), .A2(new_n678), .A3(new_n618), .ZN(new_n686));
  INV_X1    g500(.A(new_n627), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n589), .A2(new_n595), .A3(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n657), .A2(new_n688), .A3(new_n385), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n689), .A3(KEYINPUT106), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n652), .B1(new_n570), .B2(new_n572), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n649), .A3(new_n624), .A4(new_n654), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n677), .A2(new_n678), .A3(new_n618), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  OAI21_X1  g511(.A(new_n540), .B1(new_n562), .B2(new_n563), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n550), .A2(new_n565), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n698), .A2(new_n565), .B1(new_n699), .B2(new_n539), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n655), .B2(new_n656), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n381), .A2(new_n703), .A3(new_n384), .A4(new_n382), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n381), .A2(new_n384), .A3(new_n382), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n702), .A2(new_n654), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT108), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n570), .A2(new_n572), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n575), .B1(new_n709), .B2(new_n701), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n706), .A2(new_n704), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n320), .A3(new_n510), .A4(new_n649), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n317), .A2(KEYINPUT32), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n313), .A2(new_n300), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(KEYINPUT42), .A3(new_n682), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n688), .B1(new_n708), .B2(new_n713), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  NAND4_X1  g538(.A1(new_n714), .A2(new_n320), .A3(new_n510), .A4(new_n628), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  NAND2_X1  g540(.A1(new_n430), .A2(new_n595), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT43), .ZN(new_n728));
  OR3_X1    g542(.A1(new_n583), .A2(new_n728), .A3(new_n619), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n711), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT110), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n560), .B(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND2_X1  g550(.A1(G469), .A2(G902), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n709), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(G469), .C1(new_n735), .C2(G902), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n743), .A3(new_n709), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n654), .A3(new_n632), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n734), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n745), .A2(new_n749), .A3(new_n654), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n749), .B1(new_n745), .B2(new_n654), .ZN(new_n751));
  INV_X1    g565(.A(new_n320), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n586), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n750), .A2(new_n751), .A3(new_n688), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n711), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  NAND3_X1  g570(.A1(new_n714), .A2(new_n649), .A3(new_n686), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n468), .B(KEYINPUT113), .Z(new_n758));
  AND2_X1   g572(.A1(new_n711), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n608), .A2(new_n627), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n320), .A2(new_n620), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n725), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n596), .B1(new_n758), .B2(new_n589), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n587), .A2(new_n763), .A3(new_n584), .A4(new_n583), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n621), .A2(new_n579), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n723), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n673), .B(new_n683), .C1(new_n662), .C2(new_n668), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n665), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n696), .A2(new_n629), .A3(new_n650), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n636), .A2(new_n383), .A3(new_n687), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n573), .A3(new_n575), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n644), .A2(new_n775), .A3(new_n619), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n644), .A2(new_n775), .A3(new_n778), .A4(new_n619), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n696), .A2(new_n629), .A3(new_n650), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n771), .A2(new_n784), .A3(KEYINPUT53), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n768), .B1(new_n661), .B2(new_n664), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n725), .A2(new_n757), .A3(new_n761), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n765), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n723), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n780), .A2(new_n783), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n785), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n715), .A2(new_n716), .B1(new_n721), .B2(new_n720), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n789), .A3(new_n765), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n780), .A3(new_n783), .A4(new_n788), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n798), .B2(new_n787), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n771), .A2(new_n784), .A3(KEYINPUT116), .A4(KEYINPUT53), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT114), .B1(new_n767), .B2(new_n770), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n803), .A3(new_n788), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n784), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n787), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n794), .B1(new_n807), .B2(KEYINPUT54), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n719), .A2(new_n682), .ZN(new_n809));
  INV_X1    g623(.A(new_n728), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n658), .A2(new_n471), .A3(new_n711), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT48), .Z(new_n813));
  NAND3_X1  g627(.A1(new_n645), .A2(new_n811), .A3(new_n510), .ZN(new_n814));
  OAI211_X1 g628(.A(G952), .B(new_n361), .C1(new_n814), .C2(new_n663), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n810), .A2(new_n679), .A3(new_n471), .A4(new_n682), .ZN(new_n816));
  INV_X1    g630(.A(new_n692), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n750), .A2(new_n751), .B1(new_n576), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n711), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n638), .A2(new_n658), .A3(new_n635), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT118), .Z(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n816), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT50), .B1(new_n821), .B2(new_n816), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n811), .A2(new_n686), .A3(new_n810), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n648), .A2(new_n430), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n824), .B(new_n825), .C1(new_n814), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT117), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n813), .B(new_n815), .C1(new_n828), .C2(KEYINPUT51), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(KEYINPUT51), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n808), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n816), .A2(new_n385), .A3(new_n657), .ZN(new_n832));
  OAI22_X1  g646(.A1(new_n831), .A2(new_n832), .B1(G952), .B2(G953), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n817), .A2(KEYINPUT49), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n727), .A2(new_n635), .A3(new_n577), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n682), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT111), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n817), .A2(KEYINPUT49), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT112), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n638), .A3(new_n645), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(new_n840), .ZN(G75));
  AOI21_X1  g655(.A(new_n310), .B1(new_n785), .B2(new_n793), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(G210), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n356), .A2(new_n365), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n363), .ZN(new_n846));
  XOR2_X1   g660(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n843), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n843), .B2(new_n844), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n361), .A2(G952), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G51));
  XOR2_X1   g666(.A(new_n737), .B(KEYINPUT57), .Z(new_n853));
  AOI21_X1  g667(.A(new_n786), .B1(new_n785), .B2(new_n793), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n794), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n567), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n842), .A2(G469), .A3(new_n735), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(G54));
  NAND4_X1  g672(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .A4(new_n425), .ZN(new_n859));
  INV_X1    g673(.A(new_n851), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n785), .A2(new_n793), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n863));
  INV_X1    g677(.A(new_n425), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n861), .A2(new_n866), .A3(new_n871), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(G60));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT59), .Z(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n794), .B2(new_n854), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n591), .A2(new_n592), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n808), .B2(new_n875), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT122), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n878), .C1(new_n808), .C2(new_n875), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n881), .B2(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT123), .Z(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT60), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n785), .B2(new_n793), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n851), .B1(new_n888), .B2(new_n616), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(KEYINPUT61), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n889), .B(new_n892), .C1(new_n507), .C2(new_n888), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(KEYINPUT61), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT125), .Z(new_n895));
  XOR2_X1   g709(.A(new_n893), .B(new_n895), .Z(G66));
  AOI21_X1  g710(.A(new_n361), .B1(new_n473), .B2(G224), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n788), .A2(new_n766), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT126), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(new_n361), .ZN(new_n900));
  INV_X1    g714(.A(G898), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n845), .B1(new_n901), .B2(G953), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n900), .B(new_n902), .ZN(G69));
  NAND3_X1  g717(.A1(new_n809), .A2(new_n383), .A3(new_n636), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n734), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n905), .A2(new_n654), .A3(new_n632), .A4(new_n745), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n796), .A2(new_n782), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n755), .A3(new_n725), .A4(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n284), .B(new_n414), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n320), .B(new_n510), .C1(new_n912), .C2(new_n763), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n633), .B(new_n913), .C1(new_n912), .C2(new_n763), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n711), .B1(new_n754), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n646), .A2(new_n782), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT62), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n747), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(G953), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n625), .B1(new_n910), .B2(new_n542), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n361), .B1(new_n909), .B2(G227), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n911), .A2(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G72));
  NAND2_X1  g736(.A1(G472), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT63), .Z(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n908), .B2(new_n899), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n639), .A2(new_n193), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n918), .B2(new_n899), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n851), .B1(new_n928), .B2(new_n641), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n641), .A2(new_n926), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n807), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(G57));
endmodule


