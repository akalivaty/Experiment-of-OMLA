

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n587), .A2(n586), .ZN(G164) );
  BUF_X2 U551 ( .A(n879), .Z(n514) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n518), .Z(n879) );
  NOR2_X1 U553 ( .A1(G164), .A2(G1384), .ZN(n618) );
  INV_X1 U554 ( .A(KEYINPUT26), .ZN(n644) );
  NAND2_X1 U555 ( .A1(G160), .A2(G40), .ZN(n617) );
  NOR2_X1 U556 ( .A1(G651), .A2(n578), .ZN(n782) );
  NOR2_X1 U557 ( .A1(n523), .A2(n522), .ZN(G160) );
  AND2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U559 ( .A1(n874), .A2(G113), .ZN(n517) );
  INV_X1 U560 ( .A(G2105), .ZN(n519) );
  AND2_X2 U561 ( .A1(n519), .A2(G2104), .ZN(n878) );
  NAND2_X1 U562 ( .A1(G101), .A2(n878), .ZN(n515) );
  XOR2_X1 U563 ( .A(KEYINPUT23), .B(n515), .Z(n516) );
  NAND2_X1 U564 ( .A1(n517), .A2(n516), .ZN(n523) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  NAND2_X1 U566 ( .A1(G137), .A2(n514), .ZN(n521) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n519), .ZN(n875) );
  NAND2_X1 U568 ( .A1(G125), .A2(n875), .ZN(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n774) );
  NAND2_X1 U571 ( .A1(G85), .A2(n774), .ZN(n525) );
  XOR2_X1 U572 ( .A(KEYINPUT0), .B(G543), .Z(n578) );
  INV_X1 U573 ( .A(G651), .ZN(n527) );
  NOR2_X1 U574 ( .A1(n578), .A2(n527), .ZN(n778) );
  NAND2_X1 U575 ( .A1(G72), .A2(n778), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT64), .B(n526), .Z(n532) );
  NOR2_X1 U578 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n528), .Z(n775) );
  NAND2_X1 U580 ( .A1(G60), .A2(n775), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G47), .A2(n782), .ZN(n529) );
  AND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(G290) );
  NAND2_X1 U584 ( .A1(G86), .A2(n774), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G61), .A2(n775), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n778), .A2(G73), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT2), .B(n535), .Z(n536) );
  NOR2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n782), .A2(G48), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(G305) );
  NAND2_X1 U592 ( .A1(G64), .A2(n775), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G52), .A2(n782), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n547) );
  NAND2_X1 U595 ( .A1(G90), .A2(n774), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G77), .A2(n778), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U598 ( .A(KEYINPUT65), .B(n544), .ZN(n545) );
  XNOR2_X1 U599 ( .A(KEYINPUT9), .B(n545), .ZN(n546) );
  NOR2_X1 U600 ( .A1(n547), .A2(n546), .ZN(G171) );
  INV_X1 U601 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U602 ( .A(KEYINPUT72), .B(KEYINPUT6), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G63), .A2(n775), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G51), .A2(n782), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n551), .B(n550), .ZN(n558) );
  NAND2_X1 U607 ( .A1(n774), .A2(G89), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G76), .A2(n778), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n555), .ZN(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT71), .B(n556), .ZN(n557) );
  NOR2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U614 ( .A(n559), .B(KEYINPUT73), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U616 ( .A1(G91), .A2(n774), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G78), .A2(n778), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G65), .A2(n775), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G53), .A2(n782), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U623 ( .A(KEYINPUT66), .B(n567), .Z(G299) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G75), .A2(n778), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G62), .A2(n775), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n774), .A2(G88), .ZN(n570) );
  XOR2_X1 U629 ( .A(KEYINPUT78), .B(n570), .Z(n571) );
  NOR2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n782), .A2(G50), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(G303) );
  INV_X1 U633 ( .A(G303), .ZN(G166) );
  NAND2_X1 U634 ( .A1(G49), .A2(n782), .ZN(n576) );
  NAND2_X1 U635 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U637 ( .A1(n775), .A2(n577), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n578), .A2(G87), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(G288) );
  XNOR2_X1 U640 ( .A(G1986), .B(G290), .ZN(n969) );
  NAND2_X1 U641 ( .A1(G102), .A2(n878), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G138), .A2(n514), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U644 ( .A(KEYINPUT82), .B(n583), .ZN(n587) );
  NAND2_X1 U645 ( .A1(G114), .A2(n874), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G126), .A2(n875), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U648 ( .A1(n618), .A2(n617), .ZN(n719) );
  NAND2_X1 U649 ( .A1(n969), .A2(n719), .ZN(n734) );
  INV_X1 U650 ( .A(n734), .ZN(n709) );
  NAND2_X1 U651 ( .A1(G95), .A2(n878), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G131), .A2(n514), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n875), .A2(G119), .ZN(n590) );
  XOR2_X1 U655 ( .A(KEYINPUT84), .B(n590), .Z(n591) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n874), .A2(G107), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n868) );
  AND2_X1 U659 ( .A1(n868), .A2(G1991), .ZN(n603) );
  NAND2_X1 U660 ( .A1(G117), .A2(n874), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G129), .A2(n875), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n878), .A2(G105), .ZN(n597) );
  XOR2_X1 U664 ( .A(KEYINPUT38), .B(n597), .Z(n598) );
  NOR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U666 ( .A1(n514), .A2(G141), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n869) );
  AND2_X1 U668 ( .A1(n869), .A2(G1996), .ZN(n602) );
  NOR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n922) );
  INV_X1 U670 ( .A(n719), .ZN(n604) );
  NOR2_X1 U671 ( .A1(n922), .A2(n604), .ZN(n713) );
  XOR2_X1 U672 ( .A(KEYINPUT85), .B(n713), .Z(n616) );
  XNOR2_X1 U673 ( .A(KEYINPUT37), .B(G2067), .ZN(n710) );
  NAND2_X1 U674 ( .A1(G104), .A2(n878), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G140), .A2(n514), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U677 ( .A(KEYINPUT34), .B(n607), .ZN(n612) );
  NAND2_X1 U678 ( .A1(G116), .A2(n874), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G128), .A2(n875), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U681 ( .A(n610), .B(KEYINPUT35), .Z(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT36), .B(n613), .Z(n614) );
  XNOR2_X1 U684 ( .A(KEYINPUT83), .B(n614), .ZN(n889) );
  NOR2_X1 U685 ( .A1(n710), .A2(n889), .ZN(n913) );
  NAND2_X1 U686 ( .A1(n719), .A2(n913), .ZN(n716) );
  INV_X1 U687 ( .A(n716), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n732) );
  INV_X1 U689 ( .A(n732), .ZN(n707) );
  XOR2_X1 U690 ( .A(KEYINPUT86), .B(n617), .Z(n619) );
  NAND2_X2 U691 ( .A1(n619), .A2(n618), .ZN(n681) );
  NAND2_X1 U692 ( .A1(G8), .A2(n681), .ZN(n737) );
  NOR2_X1 U693 ( .A1(G1981), .A2(G305), .ZN(n620) );
  XOR2_X1 U694 ( .A(n620), .B(KEYINPUT24), .Z(n621) );
  NOR2_X1 U695 ( .A1(n737), .A2(n621), .ZN(n705) );
  XOR2_X1 U696 ( .A(G2078), .B(KEYINPUT88), .Z(n622) );
  XNOR2_X1 U697 ( .A(KEYINPUT25), .B(n622), .ZN(n995) );
  NOR2_X1 U698 ( .A1(n681), .A2(n995), .ZN(n624) );
  INV_X1 U699 ( .A(n681), .ZN(n664) );
  NOR2_X1 U700 ( .A1(n664), .A2(G1961), .ZN(n623) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n675) );
  AND2_X1 U702 ( .A1(G301), .A2(n675), .ZN(n631) );
  NOR2_X1 U703 ( .A1(n681), .A2(G2084), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT87), .B(n625), .Z(n692) );
  NOR2_X1 U705 ( .A1(G1966), .A2(n737), .ZN(n694) );
  NOR2_X1 U706 ( .A1(n692), .A2(n694), .ZN(n626) );
  XNOR2_X1 U707 ( .A(n626), .B(KEYINPUT90), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n627), .A2(G8), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n628), .B(KEYINPUT30), .ZN(n629) );
  NOR2_X1 U710 ( .A1(G168), .A2(n629), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(KEYINPUT31), .ZN(n679) );
  XNOR2_X1 U713 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G81), .A2(n774), .ZN(n633) );
  XNOR2_X1 U715 ( .A(n633), .B(KEYINPUT12), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT68), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G68), .A2(n778), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n638), .B(n637), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n775), .A2(G56), .ZN(n639) );
  XOR2_X1 U721 ( .A(KEYINPUT14), .B(n639), .Z(n640) );
  NOR2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n782), .A2(G43), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n980) );
  INV_X1 U725 ( .A(G1996), .ZN(n990) );
  NOR2_X1 U726 ( .A1(n681), .A2(n990), .ZN(n645) );
  XNOR2_X1 U727 ( .A(n645), .B(n644), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n681), .A2(G1341), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U730 ( .A1(n980), .A2(n648), .ZN(n659) );
  NAND2_X1 U731 ( .A1(G92), .A2(n774), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G79), .A2(n778), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G66), .A2(n775), .ZN(n652) );
  NAND2_X1 U735 ( .A1(G54), .A2(n782), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U738 ( .A(KEYINPUT15), .B(n655), .Z(n963) );
  INV_X1 U739 ( .A(n963), .ZN(n749) );
  NOR2_X1 U740 ( .A1(n664), .A2(G1348), .ZN(n657) );
  NOR2_X1 U741 ( .A1(G2067), .A2(n681), .ZN(n656) );
  NOR2_X1 U742 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n749), .A2(n660), .ZN(n658) );
  NAND2_X1 U744 ( .A1(n659), .A2(n658), .ZN(n662) );
  OR2_X1 U745 ( .A1(n660), .A2(n749), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U747 ( .A(KEYINPUT89), .B(n663), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n664), .A2(G2072), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n665), .B(KEYINPUT27), .ZN(n667) );
  AND2_X1 U750 ( .A1(G1956), .A2(n681), .ZN(n666) );
  NOR2_X1 U751 ( .A1(n667), .A2(n666), .ZN(n670) );
  INV_X1 U752 ( .A(G299), .ZN(n786) );
  NAND2_X1 U753 ( .A1(n670), .A2(n786), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U755 ( .A1(n670), .A2(n786), .ZN(n671) );
  XOR2_X1 U756 ( .A(n671), .B(KEYINPUT28), .Z(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U758 ( .A(n674), .B(KEYINPUT29), .ZN(n677) );
  NOR2_X1 U759 ( .A1(G301), .A2(n675), .ZN(n676) );
  NOR2_X1 U760 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n693) );
  INV_X1 U762 ( .A(n693), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n680), .A2(G286), .ZN(n689) );
  INV_X1 U764 ( .A(G8), .ZN(n687) );
  NOR2_X1 U765 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U766 ( .A(KEYINPUT91), .B(n682), .ZN(n685) );
  NOR2_X1 U767 ( .A1(G1971), .A2(n737), .ZN(n683) );
  NOR2_X1 U768 ( .A1(G166), .A2(n683), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n685), .A2(n684), .ZN(n686) );
  OR2_X1 U770 ( .A1(n687), .A2(n686), .ZN(n688) );
  AND2_X1 U771 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U772 ( .A(KEYINPUT92), .B(KEYINPUT32), .ZN(n690) );
  XNOR2_X1 U773 ( .A(n691), .B(n690), .ZN(n698) );
  NAND2_X1 U774 ( .A1(n692), .A2(G8), .ZN(n696) );
  NOR2_X1 U775 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U776 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U777 ( .A1(n698), .A2(n697), .ZN(n724) );
  NOR2_X1 U778 ( .A1(G2090), .A2(G303), .ZN(n699) );
  XOR2_X1 U779 ( .A(KEYINPUT95), .B(n699), .Z(n700) );
  NAND2_X1 U780 ( .A1(G8), .A2(n700), .ZN(n701) );
  NAND2_X1 U781 ( .A1(n724), .A2(n701), .ZN(n702) );
  NAND2_X1 U782 ( .A1(n702), .A2(n737), .ZN(n703) );
  XOR2_X1 U783 ( .A(KEYINPUT96), .B(n703), .Z(n704) );
  NOR2_X1 U784 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U785 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U786 ( .A1(n709), .A2(n708), .ZN(n722) );
  NAND2_X1 U787 ( .A1(n710), .A2(n889), .ZN(n910) );
  NOR2_X1 U788 ( .A1(G1996), .A2(n869), .ZN(n919) );
  NOR2_X1 U789 ( .A1(G1991), .A2(n868), .ZN(n915) );
  NOR2_X1 U790 ( .A1(G1986), .A2(G290), .ZN(n711) );
  NOR2_X1 U791 ( .A1(n915), .A2(n711), .ZN(n712) );
  NOR2_X1 U792 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U793 ( .A1(n919), .A2(n714), .ZN(n715) );
  XNOR2_X1 U794 ( .A(KEYINPUT39), .B(n715), .ZN(n717) );
  NAND2_X1 U795 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U796 ( .A1(n910), .A2(n718), .ZN(n720) );
  AND2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n744) );
  NOR2_X1 U799 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U800 ( .A1(G1971), .A2(G303), .ZN(n723) );
  NOR2_X1 U801 ( .A1(n965), .A2(n723), .ZN(n725) );
  NAND2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U803 ( .A(KEYINPUT93), .B(n726), .Z(n727) );
  NAND2_X1 U804 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NAND2_X1 U805 ( .A1(n727), .A2(n966), .ZN(n728) );
  XNOR2_X1 U806 ( .A(n728), .B(KEYINPUT94), .ZN(n739) );
  NAND2_X1 U807 ( .A1(n965), .A2(KEYINPUT33), .ZN(n729) );
  NOR2_X1 U808 ( .A1(n729), .A2(n737), .ZN(n731) );
  XOR2_X1 U809 ( .A(G1981), .B(G305), .Z(n960) );
  INV_X1 U810 ( .A(n960), .ZN(n730) );
  NOR2_X1 U811 ( .A1(n731), .A2(n730), .ZN(n733) );
  AND2_X1 U812 ( .A1(n733), .A2(n732), .ZN(n735) );
  AND2_X1 U813 ( .A1(n735), .A2(n734), .ZN(n740) );
  INV_X1 U814 ( .A(n740), .ZN(n736) );
  OR2_X1 U815 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U816 ( .A1(n739), .A2(n738), .ZN(n742) );
  AND2_X1 U817 ( .A1(n740), .A2(KEYINPUT33), .ZN(n741) );
  NOR2_X1 U818 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U820 ( .A(n745), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U821 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U822 ( .A(G57), .ZN(G237) );
  INV_X1 U823 ( .A(G132), .ZN(G219) );
  NAND2_X1 U824 ( .A1(G7), .A2(G661), .ZN(n747) );
  XNOR2_X1 U825 ( .A(n747), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U826 ( .A(G223), .ZN(n813) );
  NAND2_X1 U827 ( .A1(n813), .A2(G567), .ZN(n748) );
  XOR2_X1 U828 ( .A(KEYINPUT11), .B(n748), .Z(G234) );
  INV_X1 U829 ( .A(G860), .ZN(n773) );
  OR2_X1 U830 ( .A1(n980), .A2(n773), .ZN(G153) );
  INV_X1 U831 ( .A(G868), .ZN(n794) );
  NAND2_X1 U832 ( .A1(n749), .A2(n794), .ZN(n750) );
  XNOR2_X1 U833 ( .A(n750), .B(KEYINPUT70), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G868), .A2(G301), .ZN(n751) );
  NAND2_X1 U835 ( .A1(n752), .A2(n751), .ZN(G284) );
  NOR2_X1 U836 ( .A1(G299), .A2(G868), .ZN(n754) );
  NOR2_X1 U837 ( .A1(G286), .A2(n794), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n754), .A2(n753), .ZN(G297) );
  NAND2_X1 U839 ( .A1(n773), .A2(G559), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n755), .A2(n963), .ZN(n756) );
  XNOR2_X1 U841 ( .A(n756), .B(KEYINPUT75), .ZN(n758) );
  XOR2_X1 U842 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n757) );
  XNOR2_X1 U843 ( .A(n758), .B(n757), .ZN(G148) );
  NOR2_X1 U844 ( .A1(G868), .A2(n980), .ZN(n761) );
  NAND2_X1 U845 ( .A1(G868), .A2(n963), .ZN(n759) );
  NOR2_X1 U846 ( .A1(G559), .A2(n759), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n761), .A2(n760), .ZN(G282) );
  NAND2_X1 U848 ( .A1(G99), .A2(n878), .ZN(n763) );
  NAND2_X1 U849 ( .A1(G111), .A2(n874), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U851 ( .A(KEYINPUT76), .B(n764), .ZN(n769) );
  NAND2_X1 U852 ( .A1(G123), .A2(n875), .ZN(n765) );
  XNOR2_X1 U853 ( .A(n765), .B(KEYINPUT18), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n514), .A2(G135), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n914) );
  XNOR2_X1 U857 ( .A(n914), .B(G2096), .ZN(n771) );
  INV_X1 U858 ( .A(G2100), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(G156) );
  NAND2_X1 U860 ( .A1(G559), .A2(n963), .ZN(n772) );
  XOR2_X1 U861 ( .A(n980), .B(n772), .Z(n792) );
  NAND2_X1 U862 ( .A1(n773), .A2(n792), .ZN(n785) );
  NAND2_X1 U863 ( .A1(G93), .A2(n774), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G67), .A2(n775), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G80), .A2(n778), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT77), .B(n779), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n782), .A2(G55), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n795) );
  XNOR2_X1 U871 ( .A(n785), .B(n795), .ZN(G145) );
  XNOR2_X1 U872 ( .A(G166), .B(G305), .ZN(n789) );
  XNOR2_X1 U873 ( .A(G290), .B(n786), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(n795), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U876 ( .A(KEYINPUT19), .B(n790), .ZN(n791) );
  XNOR2_X1 U877 ( .A(n791), .B(G288), .ZN(n894) );
  XNOR2_X1 U878 ( .A(n792), .B(n894), .ZN(n793) );
  NOR2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n797) );
  NOR2_X1 U880 ( .A1(G868), .A2(n795), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(G295) );
  NAND2_X1 U882 ( .A1(G2078), .A2(G2084), .ZN(n798) );
  XOR2_X1 U883 ( .A(KEYINPUT20), .B(n798), .Z(n799) );
  NAND2_X1 U884 ( .A1(G2090), .A2(n799), .ZN(n800) );
  XNOR2_X1 U885 ( .A(KEYINPUT21), .B(n800), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n801), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U887 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U888 ( .A(KEYINPUT67), .B(G82), .ZN(G220) );
  NOR2_X1 U889 ( .A1(G219), .A2(G220), .ZN(n802) );
  XOR2_X1 U890 ( .A(KEYINPUT22), .B(n802), .Z(n803) );
  NOR2_X1 U891 ( .A1(G218), .A2(n803), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G96), .A2(n804), .ZN(n818) );
  NAND2_X1 U893 ( .A1(G2106), .A2(n818), .ZN(n808) );
  NAND2_X1 U894 ( .A1(G108), .A2(G120), .ZN(n805) );
  NOR2_X1 U895 ( .A1(G237), .A2(n805), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G69), .A2(n806), .ZN(n819) );
  NAND2_X1 U897 ( .A1(G567), .A2(n819), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U899 ( .A(KEYINPUT79), .B(n809), .ZN(G319) );
  INV_X1 U900 ( .A(G319), .ZN(n898) );
  NAND2_X1 U901 ( .A1(G661), .A2(G483), .ZN(n810) );
  XNOR2_X1 U902 ( .A(KEYINPUT80), .B(n810), .ZN(n811) );
  NOR2_X1 U903 ( .A1(n898), .A2(n811), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n815), .A2(G36), .ZN(n812) );
  XOR2_X1 U905 ( .A(KEYINPUT81), .B(n812), .Z(G176) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U911 ( .A(KEYINPUT99), .B(n817), .Z(G188) );
  XOR2_X1 U912 ( .A(G120), .B(KEYINPUT100), .Z(G236) );
  INV_X1 U914 ( .A(G108), .ZN(G238) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  NOR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  XOR2_X1 U918 ( .A(G2454), .B(G2435), .Z(n821) );
  XNOR2_X1 U919 ( .A(G2438), .B(G2427), .ZN(n820) );
  XNOR2_X1 U920 ( .A(n821), .B(n820), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT97), .B(G2446), .Z(n823) );
  XNOR2_X1 U922 ( .A(G2443), .B(G2430), .ZN(n822) );
  XNOR2_X1 U923 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U924 ( .A(n824), .B(G2451), .Z(n826) );
  XNOR2_X1 U925 ( .A(G1348), .B(G1341), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U928 ( .A1(n829), .A2(G14), .ZN(n830) );
  XOR2_X1 U929 ( .A(KEYINPUT98), .B(n830), .Z(G401) );
  XOR2_X1 U930 ( .A(G2100), .B(G2096), .Z(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2072), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2090), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1966), .B(G1956), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1981), .B(G1976), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U942 ( .A(G1971), .B(G1986), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U946 ( .A(KEYINPUT101), .B(G2474), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U948 ( .A(G1961), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n875), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n849), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U952 ( .A1(G100), .A2(n878), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n850), .B(KEYINPUT102), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G136), .A2(n514), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G112), .A2(n874), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U958 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G103), .A2(n878), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G139), .A2(n514), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G115), .A2(n874), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G127), .A2(n875), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U967 ( .A(KEYINPUT104), .B(n864), .ZN(n905) );
  XOR2_X1 U968 ( .A(KEYINPUT48), .B(KEYINPUT105), .Z(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT103), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n867), .B(G162), .Z(n871) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(G164), .B(n872), .Z(n873) );
  XNOR2_X1 U975 ( .A(n905), .B(n873), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G118), .A2(n874), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G130), .A2(n875), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G106), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G142), .A2(n514), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U985 ( .A(G160), .B(n914), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U988 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U989 ( .A(n980), .B(KEYINPUT106), .ZN(n893) );
  XNOR2_X1 U990 ( .A(G171), .B(n963), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n894), .B(G286), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G397) );
  OR2_X1 U995 ( .A1(G401), .A2(n898), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT49), .B(n899), .Z(n900) );
  XNOR2_X1 U998 ( .A(n900), .B(KEYINPUT107), .ZN(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G69), .ZN(G235) );
  INV_X1 U1004 ( .A(KEYINPUT55), .ZN(n931) );
  XNOR2_X1 U1005 ( .A(G2072), .B(KEYINPUT109), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1007 ( .A(G164), .B(G2078), .Z(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(KEYINPUT50), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n927) );
  XNOR2_X1 U1012 ( .A(G160), .B(G2084), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n925) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n920), .Z(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT108), .B(n921), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT110), .B(n928), .ZN(n929) );
  XOR2_X1 U1023 ( .A(KEYINPUT52), .B(n929), .Z(n930) );
  NAND2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(n932), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1026 ( .A(G1986), .B(G24), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1976), .B(KEYINPUT124), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(n933), .B(G23), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(G22), .B(G1971), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT125), .B(n936), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT58), .B(n939), .Z(n956) );
  XNOR2_X1 U1034 ( .A(G1348), .B(KEYINPUT59), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(G4), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(G1981), .B(G6), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(G1341), .B(G19), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1040 ( .A(KEYINPUT121), .B(G1956), .Z(n945) );
  XNOR2_X1 U1041 ( .A(G20), .B(n945), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT60), .B(n948), .Z(n950) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G21), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT122), .B(n951), .Z(n953) );
  XNOR2_X1 U1047 ( .A(G1961), .B(G5), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT123), .B(n954), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT126), .ZN(n958) );
  XOR2_X1 U1052 ( .A(n958), .B(KEYINPUT61), .Z(n1018) );
  INV_X1 U1053 ( .A(KEYINPUT120), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n1018), .A2(n959), .ZN(n988) );
  XNOR2_X1 U1055 ( .A(G168), .B(G1966), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT57), .B(n962), .Z(n986) );
  XNOR2_X1 U1058 ( .A(G1348), .B(n963), .ZN(n979) );
  XNOR2_X1 U1059 ( .A(G301), .B(G1961), .ZN(n977) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G166), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n964), .B(KEYINPUT116), .ZN(n971) );
  INV_X1 U1062 ( .A(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1066 ( .A(G1956), .B(G299), .Z(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT115), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(KEYINPUT117), .B(n975), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G1341), .B(n980), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT118), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT119), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n1016) );
  NOR2_X1 U1077 ( .A1(KEYINPUT56), .A2(n1016), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(G16), .A2(n989), .ZN(n1015) );
  XOR2_X1 U1080 ( .A(G2090), .B(G35), .Z(n1006) );
  XNOR2_X1 U1081 ( .A(G32), .B(n990), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G2067), .B(G26), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G2072), .B(G33), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G27), .B(n995), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT112), .B(n996), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(G1991), .B(G25), .Z(n999) );
  NAND2_X1 U1090 ( .A1(n999), .A2(G28), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT111), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(KEYINPUT113), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(n1004), .B(KEYINPUT53), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G34), .B(G2084), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT54), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT55), .B(n1010), .Z(n1011) );
  NOR2_X1 U1100 ( .A1(G29), .A2(n1011), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT114), .B(n1012), .Z(n1013) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1023) );
  INV_X1 U1104 ( .A(n1016), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(KEYINPUT56), .ZN(n1020) );
  OR2_X1 U1106 ( .A1(KEYINPUT120), .A2(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(G16), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

