//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  AOI21_X1  g004(.A(G101), .B1(new_n189), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n191), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT77), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n191), .A3(new_n194), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G128), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n202), .B1(new_n200), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n189), .A2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n189), .A2(KEYINPUT78), .A3(G107), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n210), .B(new_n211), .C1(new_n189), .C2(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G101), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n199), .A2(new_n207), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT10), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT66), .B1(new_n217), .B2(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n204), .A3(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(KEYINPUT0), .B2(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n222), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n190), .A2(new_n194), .A3(new_n208), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n200), .A2(KEYINPUT0), .A3(G128), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n233), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n234), .B2(G101), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n199), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G137), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n244), .B2(G137), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n246), .A2(new_n247), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n250), .A2(new_n243), .A3(new_n248), .A4(new_n245), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n243), .A3(new_n245), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n251), .A2(new_n253), .B1(G131), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n217), .A2(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(G128), .B1(new_n256), .B2(new_n201), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n222), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n202), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n199), .A2(new_n259), .A3(KEYINPUT10), .A4(new_n213), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n216), .A2(new_n241), .A3(new_n255), .A4(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT70), .A2(G953), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT70), .A2(G953), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G227), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT76), .ZN(new_n266));
  XOR2_X1   g080(.A(G110), .B(G140), .Z(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n254), .A2(G131), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n198), .A2(new_n196), .B1(new_n212), .B2(G101), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(new_n259), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n199), .A2(new_n213), .A3(new_n207), .ZN(new_n276));
  OAI211_X1 g090(.A(KEYINPUT12), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n269), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n216), .A2(new_n241), .A3(new_n260), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n273), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n268), .B1(new_n283), .B2(new_n261), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n268), .A3(new_n261), .ZN(new_n286));
  INV_X1    g100(.A(new_n261), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n277), .B2(new_n280), .ZN(new_n288));
  OAI211_X1 g102(.A(G469), .B(new_n286), .C1(new_n288), .C2(new_n268), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n187), .A2(new_n188), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  OAI21_X1  g107(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G119), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G116), .ZN(new_n297));
  INV_X1    g111(.A(G116), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n296), .A3(G116), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(KEYINPUT80), .ZN(new_n305));
  INV_X1    g119(.A(G113), .ZN(new_n306));
  XNOR2_X1  g120(.A(G116), .B(G119), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(KEYINPUT5), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n302), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n274), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G122), .ZN(new_n311));
  INV_X1    g125(.A(new_n240), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(new_n307), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n313), .B1(new_n318), .B2(new_n302), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n300), .A2(new_n301), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n307), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT68), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n322), .A3(new_n236), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n258), .A2(new_n325), .A3(new_n202), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n233), .B2(new_n237), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT7), .ZN(new_n329));
  INV_X1    g143(.A(G224), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n327), .A2(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n327), .A2(new_n328), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n331), .A2(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n324), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n311), .B(KEYINPUT8), .ZN(new_n337));
  INV_X1    g151(.A(new_n310), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n274), .A2(new_n309), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n310), .B1(new_n312), .B2(new_n323), .ZN(new_n342));
  INV_X1    g156(.A(new_n311), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n324), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n333), .B(new_n331), .Z(new_n346));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n347), .A3(new_n343), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(G210), .B1(G237), .B2(G902), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n341), .A2(new_n349), .A3(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(G214), .B1(G237), .B2(G902), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n295), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n188), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT22), .B(G137), .Z(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT75), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n325), .A2(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n374), .B2(new_n369), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n204), .ZN(new_n376));
  OAI211_X1 g190(.A(G146), .B(new_n371), .C1(new_n374), .C2(new_n369), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(KEYINPUT72), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n379), .A3(new_n204), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n296), .B2(G128), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n382), .B(new_n383), .C1(G119), .C2(new_n203), .ZN(new_n384));
  XNOR2_X1  g198(.A(G119), .B(G128), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT24), .B(G110), .Z(new_n386));
  AOI22_X1  g200(.A1(new_n384), .A2(G110), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n380), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n372), .A2(new_n373), .A3(new_n204), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT73), .ZN(new_n390));
  OAI22_X1  g204(.A1(new_n384), .A2(G110), .B1(new_n385), .B2(new_n386), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n377), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n388), .A2(KEYINPUT74), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT74), .B1(new_n388), .B2(new_n392), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n368), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n367), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT25), .B1(new_n398), .B2(new_n188), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n400));
  AOI211_X1 g214(.A(new_n400), .B(G902), .C1(new_n395), .C2(new_n397), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n363), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n363), .A2(G902), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n406));
  INV_X1    g220(.A(G237), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n264), .A2(G210), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT27), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G101), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n233), .A2(new_n237), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n251), .A2(new_n253), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n242), .A2(G134), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n248), .B1(new_n415), .B2(new_n245), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n258), .B2(new_n202), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n273), .A2(new_n413), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT68), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT68), .B1(new_n320), .B2(new_n321), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n322), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT28), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n418), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n420), .A2(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n411), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n417), .A2(new_n414), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n434), .B(new_n435), .C1(new_n255), .C2(new_n412), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n273), .A2(new_n413), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n438), .B2(new_n434), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n431), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n425), .A3(new_n411), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT31), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n418), .A2(new_n424), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n417), .A2(new_n414), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n412), .B1(new_n414), .B2(new_n270), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT30), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n436), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n448), .B2(new_n431), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT31), .A3(new_n411), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n433), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G472), .A2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n406), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT32), .ZN(new_n455));
  INV_X1    g269(.A(new_n428), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n427), .B1(new_n418), .B2(new_n424), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n432), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n411), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT31), .B1(new_n449), .B2(new_n411), .ZN(new_n461));
  INV_X1    g275(.A(new_n431), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n447), .B2(new_n436), .ZN(new_n463));
  NOR4_X1   g277(.A1(new_n463), .A2(new_n459), .A3(new_n444), .A4(new_n442), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n460), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(KEYINPUT71), .A3(new_n452), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n454), .A2(new_n455), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n443), .A2(new_n450), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n453), .B1(new_n468), .B2(new_n460), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n418), .A2(new_n424), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n426), .B2(new_n428), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n411), .A2(KEYINPUT29), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n444), .A2(new_n411), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n458), .A2(new_n411), .B1(new_n440), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n475), .B2(KEYINPUT29), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n469), .A2(KEYINPUT32), .B1(new_n476), .B2(G472), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n405), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G952), .ZN(new_n479));
  AOI211_X1 g293(.A(G953), .B(new_n479), .C1(G234), .C2(G237), .ZN(new_n480));
  INV_X1    g294(.A(new_n264), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT87), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n293), .A2(new_n362), .A3(G953), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n217), .A2(G128), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n203), .A2(G143), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G134), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n244), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G122), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G116), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n193), .B1(new_n498), .B2(KEYINPUT14), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n298), .A2(G122), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(G116), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n501), .A3(new_n193), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n496), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n495), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G107), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n509), .B2(new_n505), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n217), .A2(KEYINPUT13), .A3(G128), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT83), .A3(new_n492), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT13), .B1(new_n217), .B2(G128), .ZN(new_n513));
  OAI221_X1 g327(.A(G134), .B1(KEYINPUT83), .B2(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n506), .A2(KEYINPUT84), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT84), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n496), .A2(new_n504), .A3(new_n516), .A4(new_n505), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n490), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n244), .B1(new_n491), .B2(new_n492), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n505), .B1(new_n507), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n504), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT84), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n510), .A2(new_n514), .ZN(new_n523));
  AND4_X1   g337(.A1(new_n517), .A2(new_n522), .A3(new_n523), .A4(new_n490), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n188), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n523), .A3(new_n517), .ZN(new_n528));
  INV_X1    g342(.A(new_n490), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n515), .A2(new_n517), .A3(new_n490), .ZN(new_n531));
  AOI21_X1  g345(.A(G902), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT85), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n489), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n488), .B1(new_n525), .B2(new_n526), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT86), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n532), .A2(KEYINPUT85), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n526), .B(G902), .C1(new_n530), .C2(new_n531), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n488), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  INV_X1    g354(.A(new_n535), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n486), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  XNOR2_X1  g358(.A(G113), .B(G122), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n189), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n372), .A2(new_n373), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n390), .B1(new_n204), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g362(.A1(KEYINPUT70), .A2(G953), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT70), .A2(G953), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(G214), .A3(new_n407), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n217), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n264), .A2(G143), .A3(G214), .A4(new_n407), .ZN(new_n553));
  NAND2_X1  g367(.A1(KEYINPUT18), .A2(G131), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT18), .A3(G131), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n548), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n248), .B1(new_n552), .B2(new_n553), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n559), .A2(KEYINPUT82), .A3(KEYINPUT17), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT82), .B1(new_n559), .B2(KEYINPUT17), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(G131), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n552), .A2(new_n553), .A3(new_n248), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n378), .A2(new_n380), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n546), .B(new_n558), .C1(new_n562), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(new_n565), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n374), .B(KEYINPUT19), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(G146), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n377), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n558), .ZN(new_n574));
  INV_X1    g388(.A(new_n546), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n544), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n578), .ZN(new_n580));
  AOI211_X1 g394(.A(KEYINPUT20), .B(new_n580), .C1(new_n569), .C2(new_n576), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n558), .B1(new_n562), .B2(new_n568), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n575), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n583), .B2(new_n569), .ZN(new_n584));
  INV_X1    g398(.A(G475), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n579), .A2(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n543), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n361), .A2(new_n478), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  OAI21_X1  g404(.A(G472), .B1(new_n451), .B2(G902), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n454), .A2(new_n591), .A3(new_n466), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n355), .A2(new_n356), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n487), .A2(new_n188), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n525), .B2(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n518), .A2(new_n524), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT33), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n598), .B2(G478), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n586), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n593), .A2(new_n600), .A3(new_n486), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n405), .A2(new_n295), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n592), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NOR3_X1   g419(.A1(new_n534), .A2(KEYINPUT86), .A3(new_n535), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n569), .A2(new_n576), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT20), .B1(new_n609), .B2(new_n580), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n577), .A2(new_n544), .A3(new_n578), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT88), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT88), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n579), .B2(new_n581), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n584), .A2(new_n585), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n486), .B(KEYINPUT89), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n608), .A2(new_n615), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT90), .ZN(new_n620));
  INV_X1    g434(.A(new_n356), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n353), .B2(new_n354), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n536), .A2(new_n542), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n616), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT90), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n615), .A4(new_n618), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n620), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n592), .A2(new_n602), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT35), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  OR2_X1    g445(.A1(new_n393), .A2(new_n394), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n403), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n402), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n361), .A2(new_n588), .A3(new_n592), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(new_n637), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n641), .A2(new_n593), .A3(new_n295), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n467), .A2(new_n477), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n480), .B1(new_n484), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n624), .A2(new_n615), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n203), .ZN(G30));
  XOR2_X1   g464(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n355), .B(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n586), .A3(new_n608), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT92), .B(KEYINPUT39), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n646), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n292), .A2(new_n294), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n653), .A2(new_n657), .A3(new_n621), .A4(new_n637), .ZN(new_n658));
  INV_X1    g472(.A(new_n470), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n474), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n411), .B1(new_n463), .B2(new_n444), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n469), .A2(KEYINPUT32), .B1(G472), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n467), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n658), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT93), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  NAND3_X1  g482(.A1(new_n586), .A2(new_n599), .A3(new_n647), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT94), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n644), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n204), .ZN(G48));
  INV_X1    g486(.A(new_n405), .ZN(new_n673));
  INV_X1    g487(.A(new_n294), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n188), .B1(new_n281), .B2(new_n284), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT95), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n285), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(KEYINPUT95), .A3(G469), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n643), .A2(new_n673), .A3(new_n601), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  AOI21_X1  g497(.A(new_n593), .B1(new_n619), .B2(KEYINPUT90), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n478), .A3(new_n626), .A4(new_n680), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND2_X1  g500(.A1(new_n678), .A2(new_n679), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(new_n294), .A3(new_n622), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n543), .A2(new_n637), .A3(new_n587), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n643), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  OAI22_X1  g506(.A1(new_n461), .A2(new_n464), .B1(new_n411), .B2(new_n471), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n452), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n591), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n405), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n608), .A2(new_n622), .A3(new_n586), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n698), .A3(new_n618), .A4(new_n680), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  NAND2_X1  g514(.A1(new_n465), .A2(new_n188), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n701), .A2(G472), .B1(new_n452), .B2(new_n693), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT96), .B1(new_n702), .B2(new_n637), .ZN(new_n703));
  AND4_X1   g517(.A1(KEYINPUT96), .A2(new_n591), .A3(new_n637), .A4(new_n694), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n670), .B(new_n688), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  INV_X1    g520(.A(KEYINPUT98), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT97), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n708), .B1(new_n295), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n292), .A2(KEYINPUT97), .A3(new_n294), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n707), .A3(new_n711), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n477), .B1(KEYINPUT32), .B2(new_n469), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n673), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n718), .A3(KEYINPUT42), .A4(new_n670), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n295), .A2(new_n709), .ZN(new_n721));
  INV_X1    g535(.A(new_n708), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n707), .A2(new_n721), .A3(new_n711), .A4(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n478), .B(new_n670), .C1(new_n723), .C2(new_n712), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT99), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n724), .B2(KEYINPUT99), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT100), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n715), .A2(new_n730), .A3(new_n478), .A4(new_n670), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n725), .A3(new_n732), .A4(new_n727), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n720), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n248), .ZN(G33));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n715), .A2(new_n736), .A3(new_n478), .A4(new_n648), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n478), .B(new_n648), .C1(new_n723), .C2(new_n712), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT101), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT102), .B(G134), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G36));
  INV_X1    g556(.A(new_n268), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n280), .A2(new_n277), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(new_n287), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n745), .A2(new_n286), .ZN(new_n746));
  OAI21_X1  g560(.A(G469), .B1(new_n746), .B2(KEYINPUT45), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n747), .A2(KEYINPUT103), .B1(KEYINPUT45), .B2(new_n746), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n748), .B2(new_n749), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT46), .B(new_n291), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(new_n285), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(KEYINPUT105), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(KEYINPUT105), .A3(new_n285), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n751), .A2(new_n752), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n290), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n294), .A3(new_n655), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n587), .A2(new_n599), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n637), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(new_n592), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT107), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n722), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT106), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n762), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT108), .B(G137), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G39));
  NAND3_X1  g591(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n294), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n294), .B1(new_n755), .B2(new_n760), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n670), .A2(new_n405), .A3(new_n722), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n643), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT110), .B(G140), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G42));
  NAND2_X1  g605(.A1(new_n765), .A2(new_n480), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n405), .A3(new_n695), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n652), .A2(new_n356), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n680), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT50), .Z(new_n796));
  NAND2_X1  g610(.A1(new_n680), .A2(new_n722), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n703), .A2(new_n704), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n673), .A2(new_n480), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n664), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n586), .A2(new_n599), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n798), .A2(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n796), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n687), .A2(new_n674), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n778), .A2(new_n781), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n793), .A2(new_n722), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n798), .A2(new_n718), .ZN(new_n812));
  XOR2_X1   g626(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n586), .A3(new_n599), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n479), .B(G953), .C1(new_n793), .C2(new_n688), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n796), .A2(new_n803), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n782), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n778), .A2(KEYINPUT116), .A3(new_n781), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n805), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n818), .B1(new_n822), .B2(new_n808), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n811), .B(new_n817), .C1(new_n823), .C2(KEYINPUT51), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n539), .A2(new_n541), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n708), .A2(new_n616), .A3(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n615), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n292), .A2(new_n294), .A3(new_n647), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n643), .A3(new_n637), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n723), .A2(new_n712), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n670), .B1(new_n703), .B2(new_n704), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n737), .B2(new_n739), .ZN(new_n834));
  INV_X1    g648(.A(new_n628), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n359), .A2(new_n360), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n600), .A2(KEYINPUT112), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n600), .A2(KEYINPUT112), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n587), .A2(new_n825), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n835), .A2(new_n836), .A3(new_n618), .A4(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n841), .A2(new_n589), .A3(new_n638), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n681), .A2(new_n699), .A3(new_n691), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n643), .A2(new_n673), .A3(new_n680), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n627), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n834), .A2(new_n842), .A3(KEYINPUT53), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n734), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n642), .B(new_n643), .C1(new_n670), .C2(new_n648), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n829), .B2(new_n641), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n828), .A2(new_n637), .A3(KEYINPUT113), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n664), .B(new_n698), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n853), .A3(new_n705), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n857), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n849), .A2(new_n705), .A3(KEYINPUT52), .A4(new_n853), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n848), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n843), .B2(new_n845), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n687), .A2(new_n294), .A3(new_n622), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n689), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n283), .A2(new_n261), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n744), .A2(new_n269), .B1(new_n870), .B2(new_n268), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n187), .B1(new_n871), .B2(new_n188), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n285), .A2(new_n677), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n679), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n294), .B(new_n618), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n697), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n643), .A2(new_n869), .B1(new_n877), .B2(new_n696), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(KEYINPUT111), .A3(new_n681), .A4(new_n685), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n834), .A3(new_n842), .ZN(new_n881));
  INV_X1    g695(.A(new_n861), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n734), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n864), .B(new_n865), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n883), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n729), .A2(new_n733), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n888), .B2(new_n719), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n889), .B2(new_n863), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n891), .B2(new_n865), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n824), .A2(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n673), .A2(new_n357), .A3(new_n294), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n652), .A3(new_n763), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n687), .B(KEYINPUT49), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n664), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n264), .A2(G952), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n864), .B1(new_n883), .B2(new_n885), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G902), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n345), .A2(new_n348), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT119), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n346), .B(KEYINPUT55), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(KEYINPUT120), .A2(KEYINPUT121), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n909), .B(new_n910), .C1(KEYINPUT120), .C2(new_n903), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n903), .A2(new_n912), .A3(new_n910), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n907), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n899), .B1(new_n911), .B2(new_n914), .ZN(G51));
  AOI21_X1  g729(.A(new_n885), .B1(new_n889), .B2(new_n861), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n862), .A2(new_n734), .A3(new_n847), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT54), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n886), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n900), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n290), .B(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(KEYINPUT123), .A3(new_n871), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n902), .A2(new_n758), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n871), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n899), .B1(new_n926), .B2(new_n929), .ZN(G54));
  NAND2_X1  g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n901), .A2(new_n609), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n899), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n609), .B1(new_n901), .B2(new_n931), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(G60));
  NAND2_X1  g751(.A1(new_n919), .A2(new_n921), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n594), .B(KEYINPUT59), .ZN(new_n939));
  OR3_X1    g753(.A1(new_n938), .A2(new_n598), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n892), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n598), .B1(new_n941), .B2(new_n939), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n940), .A2(new_n933), .A3(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT60), .Z(new_n945));
  NAND4_X1  g759(.A1(new_n900), .A2(new_n635), .A3(new_n634), .A4(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n900), .A2(new_n945), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n398), .B(KEYINPUT125), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n933), .B(new_n946), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(KEYINPUT126), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT127), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G66));
  OAI21_X1  g768(.A(G953), .B1(new_n485), .B2(new_n330), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n880), .A2(new_n842), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n481), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n905), .B1(G898), .B2(new_n264), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  AOI21_X1  g773(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n762), .A2(new_n697), .A3(new_n717), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n849), .A2(new_n705), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n740), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n762), .B2(new_n774), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n961), .A2(new_n964), .A3(new_n734), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n789), .A2(new_n264), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n448), .B(new_n571), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(G900), .B2(new_n481), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n967), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n667), .A2(new_n962), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n656), .A2(new_n708), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n840), .A2(new_n478), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n775), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n789), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n970), .B1(new_n978), .B2(new_n264), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n960), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n264), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n967), .ZN(new_n982));
  INV_X1    g796(.A(new_n960), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n966), .A2(new_n968), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n985), .ZN(G72));
  NAND3_X1  g800(.A1(new_n789), .A2(new_n956), .A3(new_n977), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  AOI21_X1  g803(.A(new_n661), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n474), .A2(new_n440), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n789), .A2(new_n956), .A3(new_n965), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n989), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n661), .A2(new_n991), .A3(new_n989), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n933), .B1(new_n891), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n990), .A2(new_n993), .A3(new_n995), .ZN(G57));
endmodule


