//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n203), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n223), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT65), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n216), .ZN(new_n251));
  NAND3_X1  g0051(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT66), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT66), .A4(new_n252), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT67), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  AOI211_X1 g0063(.A(new_n263), .B(new_n260), .C1(new_n255), .C2(new_n256), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G226), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n255), .B2(new_n256), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G222), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G223), .A2(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n251), .A2(new_n248), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n268), .A2(new_n260), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n266), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G200), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n207), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G50), .ZN(new_n286));
  XOR2_X1   g0086(.A(new_n286), .B(KEYINPUT68), .Z(new_n287));
  NAND3_X1  g0087(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n216), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n277), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n294), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n204), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n291), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n289), .A2(new_n201), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT9), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n284), .B(new_n306), .C1(new_n307), .C2(new_n283), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n283), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT69), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n283), .A2(G179), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n313), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(KEYINPUT70), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n314), .A2(new_n316), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n309), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n274), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G87), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT78), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT75), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n277), .B2(KEYINPUT3), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n275), .A2(KEYINPUT75), .A3(G33), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n278), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G223), .B2(G1698), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n324), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n268), .A2(new_n260), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n257), .A2(G232), .A3(new_n261), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G169), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(G179), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n292), .ZN(new_n340));
  INV_X1    g0140(.A(new_n294), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n285), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n340), .A2(new_n342), .B1(new_n288), .B2(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(new_n291), .ZN(new_n344));
  XNOR2_X1  g0144(.A(G58), .B(G68), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n328), .A2(new_n208), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(KEYINPUT76), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n328), .B2(new_n208), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n203), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n347), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n344), .B1(new_n356), .B2(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT16), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n349), .B1(new_n269), .B2(G20), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n203), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n346), .B1(new_n361), .B2(KEYINPUT77), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n343), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT18), .B1(new_n339), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n352), .A2(new_n355), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(new_n368), .A3(new_n291), .ZN(new_n369));
  INV_X1    g0169(.A(new_n343), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n338), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n333), .B2(new_n334), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n257), .A2(G274), .A3(new_n260), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n332), .A2(new_n321), .ZN(new_n378));
  AND4_X1   g0178(.A1(G190), .A2(new_n377), .A3(new_n334), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n374), .B1(new_n365), .B2(new_n380), .ZN(new_n381));
  AND4_X1   g0181(.A1(new_n374), .A2(new_n369), .A3(new_n380), .A4(new_n370), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n366), .B(new_n373), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n265), .A2(G244), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G238), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n269), .B(new_n386), .C1(new_n226), .C2(G1698), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n274), .B1(new_n279), .B2(new_n220), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n268), .A2(new_n260), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(G169), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n295), .B1(G20), .B2(G77), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n341), .A2(new_n298), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n344), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n292), .A2(G77), .A3(new_n285), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G77), .B2(new_n288), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n390), .A2(G179), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n391), .A2(KEYINPUT71), .A3(G190), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n397), .A2(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n390), .A2(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT71), .B1(new_n391), .B2(G190), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n320), .A2(new_n384), .A3(new_n401), .A4(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n262), .A2(new_n264), .A3(new_n227), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n226), .A2(new_n270), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G97), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n411), .A2(new_n279), .B1(new_n277), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n329), .A2(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n269), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT72), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT72), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n269), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n377), .B1(new_n419), .B2(new_n274), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT13), .B1(new_n409), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n257), .A2(new_n261), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n263), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n257), .A2(KEYINPUT67), .A3(new_n261), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(G238), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(new_n418), .ZN(new_n426));
  INV_X1    g0226(.A(new_n413), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n321), .B1(new_n268), .B2(new_n260), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(G179), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n421), .A2(KEYINPUT73), .A3(new_n431), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n420), .B1(new_n265), .B2(G238), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT73), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n430), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(G169), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n434), .A2(KEYINPUT14), .A3(G169), .A4(new_n437), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n433), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n292), .A2(G68), .A3(new_n285), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n298), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n296), .B2(new_n280), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n291), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n288), .A2(G68), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT12), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(new_n451), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT74), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n454), .B2(new_n453), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n442), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n434), .A2(G200), .A3(new_n437), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n307), .B1(new_n435), .B2(new_n430), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n461), .B2(new_n421), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n408), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OR2_X1    g0266(.A1(G250), .A2(G1698), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G257), .B2(new_n270), .ZN(new_n468));
  INV_X1    g0268(.A(G294), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n328), .A2(new_n468), .B1(new_n277), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT88), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI221_X1 g0272(.A(KEYINPUT88), .B1(new_n277), .B2(new_n469), .C1(new_n328), .C2(new_n468), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n321), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT89), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n474), .B(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n207), .B(G45), .C1(new_n258), .C2(KEYINPUT5), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(KEYINPUT5), .B2(new_n258), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n255), .B2(new_n256), .ZN(new_n479));
  AOI22_X1  g0279(.A1(G264), .A2(new_n479), .B1(new_n268), .B2(new_n478), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n307), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n375), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n289), .A2(new_n220), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n485), .A2(KEYINPUT25), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(KEYINPUT25), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n291), .B(new_n289), .C1(new_n207), .C2(G33), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n486), .B(new_n487), .C1(new_n489), .C2(new_n220), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G87), .ZN(new_n492));
  NOR4_X1   g0292(.A1(new_n279), .A2(KEYINPUT22), .A3(G20), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n327), .A2(new_n278), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(new_n208), .A3(G87), .A4(new_n326), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(KEYINPUT85), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n326), .A2(new_n278), .A3(new_n327), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n208), .A4(G87), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n493), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT23), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n220), .A3(G20), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT86), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT24), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n326), .A2(new_n327), .A3(new_n208), .A4(new_n278), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT85), .B1(new_n509), .B2(new_n492), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n500), .A2(KEYINPUT22), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n493), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  INV_X1    g0314(.A(new_n507), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT87), .B1(new_n517), .B2(new_n291), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT87), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n519), .B(new_n344), .C1(new_n508), .C2(new_n516), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n484), .B(new_n491), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n288), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n488), .B2(G97), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n220), .B1(new_n412), .B2(KEYINPUT6), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G97), .A3(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G97), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n530), .A3(KEYINPUT6), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n531), .A3(G20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n298), .A2(G77), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT80), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n359), .A2(new_n360), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n540), .A2(KEYINPUT81), .A3(new_n291), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT81), .B1(new_n540), .B2(new_n291), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n523), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  INV_X1    g0344(.A(G244), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(G1698), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n269), .A2(new_n546), .B1(G33), .B2(G283), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n269), .B2(G250), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n270), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT4), .B1(new_n498), .B2(G244), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n321), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n268), .A2(new_n478), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n479), .A2(G257), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G169), .ZN(new_n555));
  INV_X1    g0355(.A(G179), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n554), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n543), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n543), .A2(KEYINPUT82), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n536), .B1(new_n532), .B2(new_n533), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n220), .B1(new_n359), .B2(new_n360), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n344), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n540), .A2(KEYINPUT81), .A3(new_n291), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n523), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n554), .A2(new_n307), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(G200), .B2(new_n554), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n559), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n528), .A2(new_n530), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT19), .B1(new_n573), .B2(new_n295), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n528), .A2(new_n530), .A3(new_n492), .A4(new_n220), .ZN(new_n575));
  NAND3_X1  g0375(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n208), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n574), .B1(new_n578), .B2(KEYINPUT83), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT83), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n580), .A3(new_n577), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n498), .A2(KEYINPUT84), .A3(new_n208), .A4(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n509), .B2(new_n203), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n291), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n394), .A2(new_n288), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n488), .A2(G87), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n259), .A2(G1), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n267), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n592), .B2(G250), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n255), .B2(new_n256), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G116), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n545), .A2(G1698), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G238), .B2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n328), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n321), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n375), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n600), .A2(new_n321), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n595), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(G190), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n488), .A2(new_n394), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n587), .A2(new_n589), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n603), .A2(new_n556), .A3(new_n595), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G169), .B1(new_n603), .B2(new_n595), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n591), .A2(new_n605), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n521), .A2(new_n558), .A3(new_n572), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n288), .A2(G116), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n488), .B2(G116), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT20), .ZN(new_n616));
  INV_X1    g0416(.A(G283), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n208), .B1(new_n277), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n573), .B2(new_n277), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n290), .A2(new_n216), .B1(G20), .B2(new_n222), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g0422(.A(KEYINPUT79), .B(G97), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(G33), .ZN(new_n624));
  OAI211_X1 g0424(.A(KEYINPUT20), .B(new_n620), .C1(new_n624), .C2(new_n618), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n615), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n221), .A2(G1698), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(G257), .B2(G1698), .ZN(new_n630));
  INV_X1    g0430(.A(G303), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n328), .A2(new_n630), .B1(new_n631), .B2(new_n269), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n479), .A2(G270), .B1(new_n321), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(G190), .A3(new_n552), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n552), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n628), .B(new_n634), .C1(new_n636), .C2(new_n375), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G179), .A3(new_n627), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT21), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n311), .B1(new_n615), .B2(new_n626), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n635), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n640), .A2(new_n635), .A3(new_n639), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n637), .B(new_n638), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n645));
  AOI211_X1 g0445(.A(KEYINPUT24), .B(new_n507), .C1(new_n511), .C2(new_n512), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n291), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n519), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n517), .A2(KEYINPUT87), .A3(new_n291), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n490), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n480), .A2(G179), .A3(new_n474), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n653));
  INV_X1    g0453(.A(new_n480), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n474), .A2(new_n475), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n474), .A2(new_n475), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n652), .B(new_n653), .C1(new_n657), .C2(new_n311), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n644), .B1(new_n650), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n466), .A2(new_n613), .A3(new_n660), .ZN(G372));
  AND2_X1   g0461(.A1(new_n366), .A2(new_n373), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n460), .A2(new_n462), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n459), .B1(new_n664), .B2(new_n401), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n381), .A2(new_n382), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n309), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n319), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n557), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n559), .B2(new_n569), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n612), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n607), .A2(new_n611), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n543), .A2(new_n557), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n612), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n638), .B1(new_n642), .B2(new_n641), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n491), .B1(new_n518), .B2(new_n520), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n658), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n674), .B(new_n678), .C1(new_n613), .C2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n670), .B1(new_n466), .B2(new_n683), .ZN(G369));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n658), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n691), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n521), .B1(new_n650), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n685), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  INV_X1    g0497(.A(new_n679), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n628), .A2(new_n693), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n679), .A2(KEYINPUT91), .A3(new_n699), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n701), .B(new_n702), .C1(new_n643), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n694), .A2(new_n685), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n698), .A2(new_n691), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n692), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n211), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G1), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n575), .A2(G116), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n214), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n682), .A2(new_n693), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT93), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n682), .A2(new_n721), .A3(new_n693), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n568), .B1(new_n567), .B2(new_n523), .ZN(new_n724));
  INV_X1    g0524(.A(new_n523), .ZN(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT82), .B(new_n725), .C1(new_n565), .C2(new_n566), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n612), .B(new_n557), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT94), .B1(new_n727), .B2(new_n673), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n672), .A2(new_n729), .A3(KEYINPUT26), .A4(new_n612), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT26), .B1(new_n676), .B2(new_n612), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n675), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT95), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n698), .B1(new_n650), .B2(new_n659), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n613), .B1(KEYINPUT96), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n681), .A2(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n735), .A2(new_n736), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n559), .A2(new_n569), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT26), .A3(new_n557), .A4(new_n612), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n731), .B1(new_n743), .B2(KEYINPUT94), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n736), .B(new_n675), .C1(new_n744), .C2(new_n730), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n691), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n723), .B1(new_n747), .B2(new_n720), .ZN(new_n748));
  INV_X1    g0548(.A(G330), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n572), .A2(new_n558), .A3(new_n612), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n643), .B1(new_n680), .B2(new_n658), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(new_n521), .A4(new_n693), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n608), .A2(new_n480), .A3(new_n474), .A4(new_n633), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT92), .B1(new_n753), .B2(new_n554), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  OAI211_X1 g0556(.A(KEYINPUT92), .B(new_n756), .C1(new_n753), .C2(new_n554), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n604), .A2(G179), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n482), .A3(new_n554), .A4(new_n635), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n760), .B2(new_n691), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n749), .B1(new_n752), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n748), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n717), .B1(new_n765), .B2(G1), .ZN(G364));
  INV_X1    g0566(.A(new_n704), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n208), .A2(G13), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n207), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n712), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n703), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n711), .A2(new_n279), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G355), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G116), .B2(new_n211), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n711), .A2(new_n498), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n259), .B2(new_n215), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n243), .A2(G45), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n208), .B1(KEYINPUT97), .B2(new_n311), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n311), .A2(KEYINPUT97), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n216), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n771), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n784), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n208), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G179), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n208), .A2(new_n556), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n307), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n798), .A2(new_n307), .A3(G200), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n201), .B1(new_n203), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n208), .B1(new_n793), .B2(G190), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT99), .Z(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G97), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n375), .A2(G179), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n792), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT98), .Z(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G107), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n208), .A2(new_n307), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n556), .A2(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n808), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n202), .A2(new_n814), .B1(new_n815), .B2(new_n492), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n792), .A2(new_n813), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n279), .B(new_n816), .C1(G77), .C2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n804), .A2(new_n807), .A3(new_n811), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n810), .A2(G283), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n279), .B1(new_n815), .B2(new_n631), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G326), .B2(new_n800), .ZN(new_n823));
  INV_X1    g0623(.A(new_n802), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT33), .B(G317), .ZN(new_n825));
  INV_X1    g0625(.A(new_n805), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n824), .A2(new_n825), .B1(new_n826), .B2(G294), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n814), .A2(new_n828), .B1(new_n817), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G329), .B2(new_n795), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n821), .A2(new_n823), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n791), .B1(new_n820), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n790), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n787), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n703), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n773), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NAND2_X1  g0638(.A1(new_n719), .A2(new_n722), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n401), .A2(new_n691), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n405), .A2(new_n406), .B1(new_n403), .B2(new_n693), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n401), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n682), .A2(new_n693), .A3(new_n842), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n764), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n771), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n844), .A2(new_n764), .A3(new_n845), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n814), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n850), .B1(new_n818), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n297), .B2(new_n802), .C1(new_n852), .C2(new_n801), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT34), .Z(new_n854));
  NAND2_X1  g0654(.A1(new_n810), .A2(G68), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n826), .A2(G58), .ZN(new_n856));
  INV_X1    g0656(.A(new_n815), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G50), .A2(new_n857), .B1(new_n795), .B2(G132), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n498), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n810), .A2(G87), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n800), .A2(G303), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n269), .B1(new_n857), .B2(G107), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G294), .A2(new_n850), .B1(new_n795), .B2(G311), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT100), .B(G283), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n802), .A2(new_n865), .B1(new_n817), .B2(new_n222), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(KEYINPUT101), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n807), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n854), .A2(new_n859), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n784), .ZN(new_n871));
  INV_X1    g0671(.A(new_n771), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n784), .A2(new_n785), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n280), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n871), .B(new_n874), .C1(new_n842), .C2(new_n786), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n849), .A2(new_n875), .ZN(G384));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n613), .A2(new_n660), .A3(new_n691), .ZN(new_n878));
  INV_X1    g0678(.A(new_n762), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n877), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n752), .A2(KEYINPUT104), .A3(new_n763), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI221_X4 g0684(.A(new_n433), .B1(new_n460), .B2(new_n462), .C1(new_n440), .C2(new_n441), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n457), .A2(new_n691), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT102), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n442), .B2(new_n463), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n463), .B(new_n886), .C1(new_n442), .C2(new_n458), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n884), .A2(new_n842), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n343), .B1(new_n896), .B2(new_n357), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n689), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n383), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n369), .A2(new_n380), .A3(new_n370), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n897), .B2(new_n689), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n897), .A2(new_n339), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n371), .A2(new_n338), .ZN(new_n904));
  INV_X1    g0704(.A(new_n689), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n371), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n904), .A2(new_n906), .A3(new_n907), .A4(new_n900), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n899), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n910));
  XOR2_X1   g0710(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n904), .A2(new_n906), .A3(new_n900), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n908), .ZN(new_n915));
  INV_X1    g0715(.A(new_n906), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n383), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n912), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n895), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n899), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n908), .A2(new_n914), .B1(new_n383), .B2(new_n916), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n920), .B(KEYINPUT105), .C1(new_n921), .C2(new_n912), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n894), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n899), .A2(new_n909), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n920), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n884), .A2(new_n842), .A3(new_n927), .A4(new_n892), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n893), .A2(new_n923), .B1(new_n928), .B2(new_n894), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n465), .A2(new_n884), .ZN(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n669), .B1(new_n748), .B2(new_n465), .ZN(new_n934));
  INV_X1    g0734(.A(new_n840), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n845), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n936), .A2(new_n892), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n927), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n459), .A2(new_n691), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n927), .A2(KEYINPUT39), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n910), .A2(new_n918), .A3(KEYINPUT39), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n663), .A2(new_n689), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n934), .B(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n933), .A2(new_n945), .B1(new_n207), .B2(new_n768), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n933), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n527), .A2(new_n531), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT35), .ZN(new_n949));
  OAI211_X1 g0749(.A(G116), .B(new_n217), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n215), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n201), .A2(G68), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n207), .B(G13), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n947), .A2(new_n952), .A3(new_n955), .ZN(G367));
  NOR2_X1   g0756(.A1(new_n239), .A2(new_n778), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n788), .B1(new_n211), .B2(new_n393), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n771), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n857), .A2(G116), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT46), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(new_n961), .B1(new_n800), .B2(G311), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .C1(new_n220), .C2(new_n805), .ZN(new_n963));
  INV_X1    g0763(.A(new_n865), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n850), .A2(G303), .B1(new_n818), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(G317), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n965), .B1(new_n966), .B2(new_n794), .C1(new_n623), .C2(new_n809), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n328), .B1(new_n802), .B2(new_n469), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n963), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n806), .A2(G68), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n800), .A2(G143), .ZN(new_n971));
  INV_X1    g0771(.A(new_n809), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n279), .B1(new_n972), .B2(G77), .ZN(new_n973));
  INV_X1    g0773(.A(G159), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(new_n973), .C1(new_n974), .C2(new_n802), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n814), .A2(new_n297), .B1(new_n817), .B2(new_n201), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n815), .A2(new_n202), .B1(new_n794), .B2(new_n852), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n969), .B1(new_n970), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n959), .B1(new_n980), .B2(new_n784), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n591), .A2(new_n693), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n612), .A2(new_n982), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n675), .A2(new_n591), .A3(new_n693), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT106), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT106), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n981), .B1(new_n988), .B2(new_n835), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n991));
  XNOR2_X1  g0791(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n742), .A2(new_n691), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n558), .A3(new_n572), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n672), .A2(new_n691), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n695), .A2(new_n708), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n999), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n558), .B1(new_n1001), .B2(new_n685), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(KEYINPUT42), .A2(new_n1000), .B1(new_n1002), .B2(new_n693), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1000), .A2(KEYINPUT42), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT109), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n995), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1010), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1013), .B(new_n994), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n706), .A2(new_n1001), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1011), .A2(new_n1014), .B1(new_n706), .B2(new_n1001), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n709), .A2(new_n999), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT45), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n709), .A2(new_n999), .A3(KEYINPUT44), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT44), .B1(new_n709), .B2(new_n999), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OR3_X1    g0824(.A1(new_n1021), .A2(new_n1024), .A3(new_n705), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n705), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n695), .A2(new_n708), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n695), .A2(new_n708), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1028), .A2(new_n704), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n704), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n765), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n712), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n770), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n989), .B1(new_n1019), .B2(new_n1036), .ZN(G387));
  AOI21_X1  g0837(.A(new_n778), .B1(new_n235), .B2(G45), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n715), .B2(new_n774), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n341), .A2(new_n201), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n259), .B1(new_n203), .B2(new_n280), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1041), .A2(new_n715), .A3(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1039), .A2(new_n1043), .B1(G107), .B2(new_n211), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n872), .B1(new_n1044), .B2(new_n788), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n815), .A2(new_n469), .B1(new_n805), .B2(new_n865), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G317), .A2(new_n850), .B1(new_n818), .B2(G303), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n829), .B2(new_n802), .C1(new_n828), .C2(new_n801), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT49), .ZN(new_n1053));
  INV_X1    g0853(.A(G326), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n328), .B1(new_n794), .B2(new_n1054), .C1(new_n222), .C2(new_n809), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1052), .B2(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n806), .A2(new_n394), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n201), .B2(new_n814), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT111), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n802), .A2(new_n294), .B1(new_n817), .B2(new_n203), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n810), .A2(G97), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n857), .A2(G77), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n795), .A2(G150), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1061), .A2(new_n498), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT110), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1060), .B(new_n1065), .C1(G159), .C2(new_n800), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1053), .A2(new_n1056), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1045), .B1(new_n1067), .B2(new_n791), .C1(new_n695), .C2(new_n835), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1032), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n770), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n765), .A2(new_n1070), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n712), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n765), .A2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(G393));
  NOR2_X1   g0875(.A1(new_n778), .A2(new_n246), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n788), .B1(new_n211), .B2(new_n623), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n771), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n269), .B1(new_n795), .B2(G322), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n857), .A2(new_n964), .B1(new_n818), .B2(G294), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n824), .A2(G303), .B1(new_n826), .B2(G116), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n811), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n800), .A2(G317), .B1(new_n850), .B2(G311), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n795), .A2(G143), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n203), .B2(new_n815), .C1(new_n294), .C2(new_n817), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n328), .B(new_n1089), .C1(G50), .C2(new_n824), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n800), .A2(G150), .B1(new_n850), .B2(G159), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n806), .A2(G77), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1090), .A2(new_n860), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1086), .A2(new_n1087), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1078), .B1(new_n1095), .B2(new_n784), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n999), .B2(new_n835), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1027), .B2(new_n769), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1072), .A2(new_n1027), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n713), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1072), .A2(new_n1027), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(G390));
  OAI21_X1  g0903(.A(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n885), .A2(KEYINPUT102), .A3(new_n886), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(G330), .B(new_n842), .C1(new_n878), .C2(new_n881), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n884), .A2(G330), .A3(new_n842), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n841), .A2(new_n401), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n840), .B1(new_n747), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n891), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n440), .A2(new_n441), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n432), .A3(new_n463), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n886), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n889), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n1107), .A3(new_n890), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n752), .A2(KEYINPUT104), .A3(new_n763), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT104), .B1(new_n752), .B2(new_n763), .ZN(new_n1122));
  OAI21_X1  g0922(.A(G330), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n842), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n936), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT115), .B1(new_n1125), .B2(new_n936), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1113), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n466), .A2(new_n1123), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n669), .B(new_n1129), .C1(new_n748), .C2(new_n465), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n941), .B1(KEYINPUT39), .B2(new_n927), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n937), .B2(new_n939), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n740), .A2(new_n1134), .A3(new_n521), .A4(new_n750), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n675), .B1(new_n744), .B2(new_n730), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(KEYINPUT95), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n693), .B(new_n1111), .C1(new_n1137), .C2(new_n745), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1106), .B1(new_n1138), .B2(new_n935), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n919), .A2(new_n922), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n459), .B2(new_n691), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1108), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1133), .B(new_n1145), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n713), .B1(new_n1131), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1128), .A2(new_n1144), .A3(new_n1130), .A4(new_n1146), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1132), .A2(new_n785), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n279), .B1(new_n492), .B2(new_n815), .C1(new_n801), .C2(new_n617), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G107), .B2(new_n824), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n814), .A2(new_n222), .B1(new_n794), .B2(new_n469), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n573), .B2(new_n818), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1153), .A2(new_n855), .A3(new_n1093), .A4(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n269), .B1(new_n809), .B2(new_n201), .C1(new_n802), .C2(new_n852), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G128), .B2(new_n800), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n806), .A2(G159), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n815), .A2(new_n297), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  INV_X1    g0961(.A(G132), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n814), .A2(new_n1162), .B1(new_n794), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n818), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n791), .B1(new_n1156), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n873), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n771), .B1(new_n1170), .B2(new_n341), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT116), .Z(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1151), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1147), .B2(new_n769), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1150), .A2(new_n1176), .ZN(G378));
  XOR2_X1   g0977(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1178));
  AND2_X1   g0978(.A1(new_n320), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n320), .A2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n310), .A2(new_n689), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR3_X1    g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n929), .B2(G330), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n928), .A2(new_n894), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n843), .B1(new_n1119), .B2(new_n890), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n923), .A2(new_n1188), .A3(new_n884), .ZN(new_n1189));
  AND4_X1   g0989(.A1(G330), .A2(new_n1187), .A3(new_n1189), .A4(new_n1185), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n944), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n1189), .A3(G330), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n929), .A2(G330), .A3(new_n1185), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n944), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n770), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n771), .B1(new_n1170), .B2(G50), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n814), .A2(new_n220), .B1(new_n817), .B2(new_n393), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n498), .A2(G41), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G283), .C2(new_n795), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1062), .B1(new_n202), .B2(new_n809), .C1(new_n412), .C2(new_n802), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G116), .B2(new_n800), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1205), .A3(new_n970), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1202), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n815), .A2(new_n1165), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1211), .A2(KEYINPUT117), .B1(new_n850), .B2(G128), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(KEYINPUT117), .B2(new_n1211), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT118), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n824), .A2(G132), .B1(new_n818), .B2(G137), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1163), .B2(new_n801), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G150), .B2(new_n806), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT59), .Z(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n972), .A2(G159), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1210), .B1(new_n1207), .B2(new_n1206), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1199), .B1(new_n1226), .B2(new_n784), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1185), .B2(new_n786), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1198), .A2(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1149), .A2(new_n1130), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n712), .B1(new_n1230), .B2(KEYINPUT57), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1149), .A2(new_n1130), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1232), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1231), .B2(new_n1233), .ZN(G375));
  NAND2_X1  g1034(.A1(new_n1125), .A2(new_n936), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT115), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n936), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1237), .A2(new_n1238), .B1(new_n1112), .B2(new_n1110), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT120), .B1(new_n1239), .B2(new_n769), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT120), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1128), .A2(new_n1241), .A3(new_n770), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1106), .A2(new_n785), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT121), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n872), .B1(new_n873), .B2(new_n203), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n279), .B1(new_n794), .B2(new_n631), .C1(new_n802), .C2(new_n222), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G294), .B2(new_n800), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n810), .A2(G77), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n814), .A2(new_n617), .B1(new_n817), .B2(new_n220), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G97), .B2(new_n857), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1057), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n806), .A2(G50), .ZN(new_n1252));
  INV_X1    g1052(.A(G128), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n814), .A2(new_n852), .B1(new_n794), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G150), .B2(new_n818), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n815), .A2(new_n974), .B1(new_n809), .B2(new_n202), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n328), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G132), .A2(new_n800), .B1(new_n824), .B2(new_n1166), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1252), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1251), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1244), .B(new_n1245), .C1(new_n791), .C2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1240), .A2(new_n1242), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1131), .A2(new_n1035), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(G381));
  OR2_X1    g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(G381), .A2(G384), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1175), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1102), .B(new_n989), .C1(new_n1036), .C2(new_n1019), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1270), .A2(G375), .A3(new_n1271), .ZN(G407));
  NAND2_X1  g1072(.A1(new_n690), .A2(G213), .ZN(new_n1273));
  OR3_X1    g1073(.A1(G375), .A2(G378), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(G213), .A3(new_n1274), .ZN(G409));
  OAI211_X1 g1075(.A(G378), .B(new_n1229), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1230), .A2(new_n1035), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1198), .A2(new_n1228), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1269), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1273), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT123), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT123), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1283), .A3(new_n1273), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n690), .A2(G213), .A3(G2897), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1129), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n693), .B1(new_n1137), .B2(new_n745), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(KEYINPUT29), .B2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n670), .B(new_n1287), .C1(new_n1290), .C2(new_n466), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1286), .A2(new_n1291), .A3(KEYINPUT60), .A4(new_n1113), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT122), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1239), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n713), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1301), .B2(new_n1263), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(G384), .A3(new_n1263), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1285), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1285), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1282), .B(new_n1284), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(G384), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1308), .B(new_n1262), .C1(new_n1296), .C2(new_n1300), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(new_n1302), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1280), .A2(new_n1273), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1280), .A2(new_n1273), .A3(new_n1310), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G393), .A2(G396), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1267), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT124), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G387), .A2(G390), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT124), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1267), .A2(new_n1316), .A3(new_n1320), .ZN(new_n1321));
  AND4_X1   g1121(.A1(new_n1271), .A2(new_n1318), .A3(new_n1319), .A4(new_n1321), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1318), .A2(new_n1321), .B1(new_n1319), .B2(new_n1271), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(KEYINPUT61), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1307), .A2(new_n1312), .A3(new_n1315), .A4(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1281), .B1(new_n1306), .B2(new_n1305), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  XOR2_X1   g1129(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1330));
  NAND2_X1  g1130(.A1(new_n1313), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT126), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1331), .A2(new_n1332), .B1(new_n1311), .B2(KEYINPUT62), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1313), .A2(KEYINPUT126), .A3(new_n1330), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1329), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1324), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1326), .B1(new_n1335), .B2(new_n1336), .ZN(G405));
  INV_X1    g1137(.A(new_n1310), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(KEYINPUT127), .ZN(new_n1339));
  OR2_X1    g1139(.A1(new_n1324), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1324), .A2(new_n1339), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  OR2_X1    g1142(.A1(new_n1338), .A2(KEYINPUT127), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1269), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1276), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1345), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(G402));
endmodule


