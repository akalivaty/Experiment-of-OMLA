//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  OAI21_X1  g005(.A(G143), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n190), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n192), .A2(new_n193), .A3(G128), .A4(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT66), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n190), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G146), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n196), .B1(new_n202), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(G137), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n215), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n208), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n211), .A2(new_n215), .A3(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n216), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n188), .A2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n206), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n229), .B2(new_n203), .ZN(new_n230));
  OR3_X1    g044(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(new_n192), .B2(new_n195), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n224), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n187), .B1(new_n220), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  OR2_X1    g054(.A1(KEYINPUT67), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT67), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n243), .B2(G116), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n241), .B2(new_n242), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n245), .B1(new_n249), .B2(new_n240), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n222), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(new_n222), .B2(new_n216), .ZN(new_n253));
  INV_X1    g067(.A(new_n233), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n230), .B2(new_n231), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n252), .A2(new_n253), .B1(new_n255), .B2(new_n235), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n208), .A2(new_n216), .A3(new_n219), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT30), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n238), .A2(new_n251), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n251), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(G101), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G953), .ZN(new_n268));
  AOI21_X1  g082(.A(G237), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G210), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n264), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n251), .B1(new_n220), .B2(new_n237), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT28), .A4(new_n260), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n273), .B(new_n274), .C1(new_n272), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n256), .A2(new_n257), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n251), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n281), .A2(KEYINPUT71), .B1(new_n284), .B2(new_n276), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n272), .A2(new_n274), .ZN(new_n286));
  AOI21_X1  g100(.A(G902), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G472), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n279), .A2(new_n272), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n259), .A2(new_n261), .A3(new_n271), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n259), .A2(new_n294), .A3(new_n261), .A4(new_n271), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n279), .A2(new_n296), .A3(new_n272), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n291), .A2(new_n293), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n289), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(G125), .A2(G140), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G125), .A2(G140), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n205), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n313), .B2(new_n305), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n309), .B1(new_n316), .B2(G146), .ZN(new_n317));
  AND2_X1   g131(.A1(KEYINPUT67), .A2(G119), .ZN(new_n318));
  NOR2_X1   g132(.A1(KEYINPUT67), .A2(G119), .ZN(new_n319));
  OAI21_X1  g133(.A(G128), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT66), .B(G128), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n320), .B(KEYINPUT23), .C1(new_n239), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n241), .A2(new_n323), .A3(new_n197), .A4(new_n242), .ZN(new_n324));
  AOI21_X1  g138(.A(G110), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(G128), .A2(new_n243), .B1(new_n201), .B2(G119), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT24), .B(G110), .Z(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n317), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT74), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n331), .B(new_n317), .C1(new_n325), .C2(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n190), .B1(new_n314), .B2(new_n315), .ZN(new_n334));
  INV_X1    g148(.A(new_n315), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n335), .B(G146), .C1(new_n308), .C2(new_n310), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT73), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n322), .A2(G110), .A3(new_n324), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n326), .A2(new_n327), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n316), .A2(new_n340), .A3(G146), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n337), .A2(new_n338), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(G137), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n266), .A2(new_n268), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(KEYINPUT75), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n333), .A2(new_n352), .A3(new_n342), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n350), .B1(new_n354), .B2(new_n349), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT72), .B(G217), .ZN(new_n356));
  INV_X1    g170(.A(G234), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G902), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n362));
  INV_X1    g176(.A(new_n350), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n333), .A2(new_n352), .A3(new_n342), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n352), .B1(new_n333), .B2(new_n342), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n366), .B2(new_n348), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n362), .B1(new_n367), .B2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n369));
  INV_X1    g183(.A(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n362), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n355), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n361), .B1(new_n373), .B2(new_n359), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n304), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n376));
  OAI21_X1  g190(.A(G116), .B1(new_n318), .B2(new_n319), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n376), .B(G113), .C1(new_n377), .C2(KEYINPUT5), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n377), .B(KEYINPUT5), .C1(G116), .C2(new_n239), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n243), .A2(new_n381), .A3(G116), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n376), .B1(new_n382), .B2(G113), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n247), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT3), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n390), .A2(new_n391), .A3(new_n393), .A4(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT80), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(G101), .C1(KEYINPUT80), .C2(new_n389), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n384), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT8), .ZN(new_n405));
  INV_X1    g219(.A(G113), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n249), .B2(new_n381), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n407), .A2(new_n379), .B1(new_n246), .B2(new_n244), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(new_n400), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n404), .A2(KEYINPUT8), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G125), .B1(new_n255), .B2(new_n235), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT1), .B1(new_n205), .B2(new_n206), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n207), .B1(new_n414), .B2(new_n321), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n206), .B1(new_n227), .B2(new_n228), .ZN(new_n416));
  NOR4_X1   g230(.A1(new_n416), .A2(KEYINPUT1), .A3(new_n197), .A4(new_n194), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n311), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n265), .A2(G224), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n419), .A2(KEYINPUT7), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n413), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n413), .B2(new_n418), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n412), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n394), .A2(KEYINPUT3), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n395), .B1(new_n396), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n393), .B1(new_n386), .B2(new_n389), .ZN(new_n427));
  OAI21_X1  g241(.A(G101), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT4), .A3(new_n398), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(G101), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n251), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n408), .A2(new_n401), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n403), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n412), .B(new_n435), .C1(new_n421), .C2(new_n422), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n424), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n404), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n442), .A3(new_n404), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n413), .A2(new_n418), .A3(new_n419), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n419), .B1(new_n413), .B2(new_n418), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n437), .A2(new_n370), .A3(new_n438), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n449));
  INV_X1    g263(.A(new_n438), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n424), .A2(new_n434), .A3(new_n436), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n370), .ZN(new_n452));
  OAI211_X1 g266(.A(KEYINPUT84), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT85), .B1(new_n450), .B2(KEYINPUT84), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n437), .A2(new_n370), .A3(new_n447), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n457), .B(KEYINPUT81), .Z(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n197), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n192), .B2(new_n195), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n398), .B(new_n400), .C1(new_n417), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n429), .B(new_n431), .C1(new_n255), .C2(new_n235), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n208), .A2(new_n401), .A3(KEYINPUT10), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n252), .A2(new_n253), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n466), .A3(new_n469), .A4(new_n467), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n346), .A2(G227), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G140), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n229), .A2(new_n203), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n227), .A2(new_n228), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n193), .B1(new_n479), .B2(G143), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n480), .B2(new_n201), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n409), .A2(new_n481), .A3(new_n196), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n463), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n469), .B1(new_n463), .B2(new_n482), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(KEYINPUT12), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n473), .A2(new_n476), .B1(new_n477), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n370), .ZN(new_n490));
  NAND2_X1  g304(.A1(G469), .A2(G902), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n483), .B2(new_n470), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n493), .B(new_n224), .C1(new_n463), .C2(new_n482), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n472), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n476), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n471), .A2(new_n472), .A3(new_n476), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(G469), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n491), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G221), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT9), .B(G234), .Z(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n370), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT78), .Z(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n201), .A2(G143), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(G134), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n197), .A2(G143), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n210), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n206), .B1(new_n198), .B2(new_n200), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n516), .A2(G134), .A3(new_n513), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n512), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT91), .B1(new_n248), .B2(G122), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n521));
  INV_X1    g335(.A(G122), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(G116), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n248), .A2(G122), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n524), .A2(G107), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(G107), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n388), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n524), .A2(G107), .A3(new_n525), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n510), .A2(new_n511), .A3(G134), .A4(new_n514), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n518), .A2(new_n528), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(KEYINPUT14), .A3(G107), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n535), .A2(new_n529), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(new_n515), .C2(new_n517), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n502), .A2(new_n265), .A3(new_n356), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n534), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n534), .B2(new_n538), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n509), .B1(new_n543), .B2(new_n370), .ZN(new_n544));
  NOR4_X1   g358(.A1(new_n541), .A2(new_n542), .A3(G902), .A4(new_n508), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g362(.A1(KEYINPUT18), .A2(G131), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT86), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(G143), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n206), .A2(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n269), .A2(new_n554), .A3(G214), .ZN(new_n555));
  INV_X1    g369(.A(new_n552), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n269), .B2(G214), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G237), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n346), .A2(G214), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n552), .ZN(new_n561));
  INV_X1    g375(.A(new_n549), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n269), .A2(new_n554), .A3(G214), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n309), .B1(G146), .B2(new_n308), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n406), .A2(new_n522), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g384(.A1(G113), .A2(G122), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n573), .A2(new_n392), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n571), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT89), .ZN(new_n577));
  AOI21_X1  g391(.A(G104), .B1(new_n577), .B2(new_n572), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT90), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n392), .B1(new_n573), .B2(new_n574), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(G104), .A3(new_n572), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G131), .B1(new_n555), .B2(new_n557), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n561), .A2(new_n214), .A3(new_n563), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n337), .A2(new_n341), .ZN(new_n589));
  OAI211_X1 g403(.A(KEYINPUT17), .B(G131), .C1(new_n555), .C2(new_n557), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n568), .B(new_n584), .C1(new_n588), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n575), .A2(new_n578), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT19), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n596), .B(new_n597), .C1(new_n306), .C2(new_n307), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n313), .A2(new_n594), .A3(new_n595), .A4(new_n305), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n336), .B1(new_n601), .B2(new_n205), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n585), .B2(new_n587), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n566), .B1(new_n558), .B2(new_n564), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n593), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n592), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(G475), .A2(G902), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n548), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n607), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT20), .B(new_n609), .C1(new_n592), .C2(new_n605), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n568), .B1(new_n588), .B2(new_n591), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n593), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n612), .B2(new_n592), .ZN(new_n613));
  INV_X1    g427(.A(G475), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n608), .A2(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n547), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G952), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(G953), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n357), .B2(new_n559), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n370), .B(new_n346), .C1(G234), .C2(G237), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT21), .B(G898), .Z(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n460), .A2(new_n506), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n375), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  NAND2_X1  g441(.A1(new_n298), .A2(new_n370), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n298), .A2(new_n300), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n506), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n632), .A2(new_n374), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n458), .B1(new_n635), .B2(new_n448), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n623), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n543), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n507), .A2(G902), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT93), .B1(new_n539), .B2(KEYINPUT94), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n534), .B2(new_n538), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n534), .A2(new_n538), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT94), .B1(new_n644), .B2(KEYINPUT93), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n645), .B2(new_n540), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n640), .B(new_n641), .C1(new_n646), .C2(new_n639), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT95), .B(G478), .ZN(new_n648));
  INV_X1    g462(.A(new_n543), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n615), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n637), .A2(new_n638), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n634), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT34), .B(G104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT96), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G6));
  AND2_X1   g471(.A1(new_n592), .A2(new_n605), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT20), .B1(new_n658), .B2(new_n609), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n606), .A2(new_n548), .A3(new_n607), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n612), .A2(new_n592), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n370), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n659), .A2(new_n660), .B1(new_n662), .B2(G475), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n623), .B(KEYINPUT97), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n547), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT98), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n615), .A2(new_n546), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n665), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n636), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n634), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NAND2_X1  g490(.A1(new_n373), .A2(new_n359), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n354), .B1(KEYINPUT36), .B2(new_n348), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT36), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n366), .A2(new_n679), .A3(new_n349), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n678), .A2(new_n680), .A3(new_n360), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n632), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n681), .B1(new_n373), .B2(new_n359), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT100), .B1(new_n686), .B2(new_n631), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n685), .A2(new_n687), .A3(new_n625), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT37), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(G110), .Z(G12));
  NAND2_X1  g504(.A1(new_n635), .A2(new_n448), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n619), .B1(new_n621), .B2(G900), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT101), .Z(new_n693));
  NOR3_X1   g507(.A1(new_n615), .A2(new_n546), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n694), .A3(new_n459), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n636), .A2(new_n697), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(new_n304), .A3(new_n633), .A4(new_n683), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  XOR2_X1   g515(.A(new_n693), .B(KEYINPUT39), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n633), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n663), .A2(new_n546), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n459), .A3(new_n686), .A4(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n456), .A2(KEYINPUT103), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n456), .A2(KEYINPUT103), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n708), .A2(KEYINPUT38), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT38), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n703), .A2(new_n704), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(G472), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n262), .A2(new_n271), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n261), .A2(new_n272), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n718), .B2(new_n283), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n715), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n630), .A2(KEYINPUT32), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n720), .B1(new_n721), .B2(new_n301), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n707), .A2(new_n714), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n206), .ZN(G45));
  INV_X1    g538(.A(new_n693), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n651), .A2(new_n615), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n651), .A2(new_n728), .A3(new_n615), .A4(new_n725), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n727), .A2(new_n636), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n683), .A2(new_n730), .A3(new_n304), .A4(new_n633), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  NAND2_X1  g546(.A1(new_n488), .A2(new_n370), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n505), .A3(new_n490), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(new_n737), .A3(new_n505), .A4(new_n490), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n375), .A2(new_n653), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  AND3_X1   g556(.A1(new_n739), .A2(new_n304), .A3(new_n374), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n673), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NAND2_X1  g559(.A1(new_n721), .A2(new_n301), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n746), .A2(new_n289), .B1(new_n677), .B2(new_n682), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n637), .A2(new_n735), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n623), .A3(new_n616), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  AND2_X1   g564(.A1(new_n636), .A2(new_n706), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n665), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT107), .B(G472), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n293), .B(new_n295), .C1(new_n285), .C2(new_n271), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n628), .A2(new_n753), .B1(new_n300), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n374), .A3(new_n739), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  AND2_X1   g571(.A1(new_n727), .A2(new_n729), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n683), .A2(new_n758), .A3(new_n748), .A4(new_n755), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT108), .B(G125), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G27));
  NAND4_X1  g575(.A1(new_n449), .A2(new_n453), .A3(new_n459), .A4(new_n455), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT110), .B1(new_n763), .B2(new_n633), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n453), .A2(new_n455), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n459), .A4(new_n449), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n633), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n375), .B(new_n758), .C1(new_n764), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n769), .B(new_n770), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(KEYINPUT42), .A3(new_n375), .A4(new_n758), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  OAI211_X1 g592(.A(new_n375), .B(new_n694), .C1(new_n764), .C2(new_n771), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n476), .B1(new_n486), .B2(new_n472), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n468), .A2(new_n470), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n477), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n498), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n491), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n788), .A2(new_n789), .A3(new_n490), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n789), .B1(new_n788), .B2(new_n490), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT46), .B1(new_n787), .B2(new_n491), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n504), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(new_n702), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n663), .A2(new_n651), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n663), .A2(new_n651), .A3(KEYINPUT43), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n683), .A2(new_n631), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n763), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n802), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n795), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  XNOR2_X1  g622(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n793), .B2(new_n504), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n788), .A2(new_n490), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n788), .A2(new_n789), .A3(new_n490), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n505), .B(new_n809), .C1(new_n815), .C2(new_n792), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n804), .A2(new_n304), .A3(new_n374), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n758), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  INV_X1    g634(.A(new_n619), .ZN(new_n821));
  INV_X1    g635(.A(new_n735), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n766), .A2(new_n821), .A3(new_n768), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n798), .B2(new_n799), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n375), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT48), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n722), .A2(new_n374), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n823), .A2(new_n827), .A3(new_n652), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n374), .A2(new_n821), .A3(new_n755), .A4(new_n800), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n748), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n618), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT120), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n734), .A2(new_n490), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n505), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n811), .A2(new_n816), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n829), .A2(new_n763), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n811), .A2(new_n816), .A3(new_n839), .A4(new_n835), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT51), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n683), .A2(new_n755), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n823), .A2(new_n827), .A3(new_n651), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n824), .A2(new_n843), .B1(new_n844), .B2(new_n663), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n735), .A2(new_n459), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n829), .B(new_n846), .C1(new_n710), .C2(new_n711), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(KEYINPUT50), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(KEYINPUT50), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n847), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n826), .B(new_n832), .C1(new_n842), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n836), .A2(new_n838), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n845), .C1(new_n851), .C2(new_n852), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n854), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n720), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n506), .B1(new_n746), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n681), .B(new_n693), .C1(new_n373), .C2(new_n359), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n751), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n700), .A2(new_n865), .A3(new_n731), .A4(new_n759), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT115), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n747), .B(new_n633), .C1(new_n699), .C2(new_n730), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n759), .A4(new_n865), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n868), .B1(new_n867), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n683), .A2(new_n758), .A3(new_n755), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n764), .B2(new_n771), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n547), .A2(new_n615), .A3(new_n693), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n763), .A2(KEYINPUT114), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n766), .A2(new_n768), .A3(new_n877), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n881), .A3(new_n633), .A4(new_n747), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n779), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n744), .A2(new_n740), .A3(new_n749), .A4(new_n756), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n668), .B1(new_n615), .B2(new_n651), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n460), .A2(new_n885), .A3(new_n664), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n634), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n688), .A3(new_n626), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n777), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT53), .B1(new_n874), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n887), .A2(new_n688), .A3(new_n626), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n740), .A2(new_n756), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n744), .A3(new_n749), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n779), .A2(new_n876), .A3(new_n882), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n866), .A2(new_n868), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n896), .A2(new_n899), .A3(new_n900), .A4(new_n777), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n891), .A2(KEYINPUT54), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n874), .B2(new_n890), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n884), .A2(KEYINPUT116), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n895), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n900), .B(new_n888), .C1(new_n884), .C2(KEYINPUT116), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n899), .A4(new_n777), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n861), .A2(new_n902), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n617), .A2(new_n265), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n861), .A2(new_n902), .A3(new_n909), .A4(KEYINPUT121), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n712), .A2(new_n504), .A3(new_n796), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n833), .B1(KEYINPUT113), .B2(KEYINPUT49), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n458), .B1(KEYINPUT113), .B2(KEYINPUT49), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n833), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n827), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n915), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n903), .A2(new_n908), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n370), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(G210), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n441), .A2(new_n443), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n446), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(KEYINPUT56), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n930), .A2(new_n931), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n930), .B2(new_n931), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n346), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  NAND2_X1  g755(.A1(new_n927), .A2(KEYINPUT54), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n942), .A2(new_n909), .B1(KEYINPUT57), .B2(new_n491), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(KEYINPUT57), .B2(new_n491), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n488), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n928), .A2(new_n370), .A3(new_n787), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(new_n658), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n658), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n940), .ZN(G60));
  INV_X1    g765(.A(new_n940), .ZN(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n507), .A2(new_n370), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n902), .B2(new_n909), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n640), .B1(new_n646), .B2(new_n639), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n952), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n942), .B2(new_n909), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n927), .A2(new_n680), .A3(new_n678), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n928), .A2(new_n963), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n952), .B(new_n965), .C1(new_n966), .C2(new_n355), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g782(.A(new_n265), .B1(new_n622), .B2(G224), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n894), .B2(new_n346), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n932), .B1(G898), .B2(new_n346), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(G69));
  NAND2_X1  g786(.A1(new_n869), .A2(new_n759), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n723), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n807), .A2(new_n819), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n804), .A2(new_n703), .ZN(new_n977));
  INV_X1    g791(.A(new_n885), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n375), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n238), .A2(new_n258), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(new_n600), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n346), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n346), .B1(G227), .B2(G900), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n795), .A2(new_n375), .A3(new_n751), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n986), .A2(new_n759), .A3(new_n869), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n976), .A2(new_n987), .A3(new_n777), .A4(new_n779), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n983), .B1(new_n988), .B2(new_n346), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(G900), .B2(new_n346), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n984), .A2(new_n985), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n985), .B1(new_n984), .B2(new_n990), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n996), .B(new_n985), .C1(new_n984), .C2(new_n990), .ZN(new_n997));
  OAI22_X1  g811(.A1(new_n992), .A2(new_n993), .B1(new_n995), .B2(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n273), .A2(new_n292), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n891), .A2(new_n901), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n988), .B2(new_n894), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n272), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n952), .B(new_n1002), .C1(new_n1004), .C2(new_n262), .ZN(new_n1005));
  INV_X1    g819(.A(new_n716), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1000), .B1(new_n980), .B2(new_n894), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(G57));
endmodule


