

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752;

  INV_X1 U375 ( .A(n370), .ZN(n633) );
  BUF_X1 U376 ( .A(n653), .Z(n354) );
  NAND2_X1 U377 ( .A1(n398), .A2(n362), .ZN(n631) );
  XNOR2_X1 U378 ( .A(n514), .B(KEYINPUT102), .ZN(n653) );
  INV_X1 U379 ( .A(n365), .ZN(n355) );
  BUF_X1 U380 ( .A(G113), .Z(n353) );
  INV_X1 U381 ( .A(KEYINPUT3), .ZN(n471) );
  NAND2_X1 U382 ( .A1(n394), .A2(n534), .ZN(n370) );
  INV_X1 U383 ( .A(n517), .ZN(n524) );
  NAND2_X1 U384 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X2 U385 ( .A(n509), .B(n355), .ZN(n517) );
  XNOR2_X2 U386 ( .A(n484), .B(KEYINPUT16), .ZN(n404) );
  XNOR2_X1 U387 ( .A(n384), .B(n500), .ZN(n581) );
  NOR2_X2 U388 ( .A1(n513), .A2(n555), .ZN(n514) );
  XNOR2_X2 U389 ( .A(n518), .B(KEYINPUT22), .ZN(n538) );
  NOR2_X2 U390 ( .A1(n581), .A2(n508), .ZN(n509) );
  XNOR2_X2 U391 ( .A(n416), .B(n415), .ZN(n484) );
  AND2_X1 U392 ( .A1(n606), .A2(n605), .ZN(n741) );
  XOR2_X1 U393 ( .A(n486), .B(n485), .Z(n487) );
  AND2_X1 U394 ( .A1(n724), .A2(n607), .ZN(n608) );
  XNOR2_X1 U395 ( .A(n372), .B(n371), .ZN(n749) );
  XNOR2_X1 U396 ( .A(n562), .B(n561), .ZN(n599) );
  NOR2_X2 U397 ( .A1(n438), .A2(n527), .ZN(n663) );
  BUF_X1 U398 ( .A(n519), .Z(n520) );
  NOR2_X1 U399 ( .A1(n552), .A2(n507), .ZN(n508) );
  XNOR2_X1 U400 ( .A(n471), .B(G101), .ZN(n416) );
  XNOR2_X1 U401 ( .A(G119), .B(G113), .ZN(n415) );
  XNOR2_X1 U402 ( .A(G902), .B(KEYINPUT15), .ZN(n461) );
  INV_X2 U403 ( .A(G953), .ZN(n742) );
  XNOR2_X2 U404 ( .A(n730), .B(n399), .ZN(n624) );
  XNOR2_X2 U405 ( .A(n404), .B(n487), .ZN(n730) );
  XNOR2_X2 U406 ( .A(n448), .B(G469), .ZN(n570) );
  NAND2_X1 U407 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U408 ( .A(n580), .ZN(n390) );
  XNOR2_X1 U409 ( .A(n684), .B(n515), .ZN(n589) );
  XNOR2_X1 U410 ( .A(n740), .B(G146), .ZN(n479) );
  XNOR2_X1 U411 ( .A(n383), .B(KEYINPUT72), .ZN(n583) );
  NOR2_X1 U412 ( .A1(n580), .A2(KEYINPUT47), .ZN(n383) );
  NAND2_X1 U413 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U414 ( .A(n752), .ZN(n378) );
  AND2_X1 U415 ( .A1(n596), .A2(n376), .ZN(n375) );
  OR2_X1 U416 ( .A1(n528), .A2(n749), .ZN(n529) );
  AND2_X1 U417 ( .A1(n541), .A2(n749), .ZN(n542) );
  XOR2_X1 U418 ( .A(G122), .B(G104), .Z(n486) );
  XNOR2_X1 U419 ( .A(G146), .B(G125), .ZN(n493) );
  XNOR2_X1 U420 ( .A(n445), .B(n444), .ZN(n740) );
  XNOR2_X1 U421 ( .A(n470), .B(KEYINPUT73), .ZN(n521) );
  XNOR2_X1 U422 ( .A(n499), .B(n498), .ZN(n695) );
  XNOR2_X1 U423 ( .A(n465), .B(n464), .ZN(n680) );
  OR2_X1 U424 ( .A1(n636), .A2(G902), .ZN(n465) );
  XNOR2_X1 U425 ( .A(n373), .B(n598), .ZN(n606) );
  XNOR2_X1 U426 ( .A(G137), .B(G140), .ZN(n457) );
  XNOR2_X1 U427 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n434) );
  XNOR2_X1 U428 ( .A(n489), .B(G134), .ZN(n445) );
  XNOR2_X1 U429 ( .A(n432), .B(n382), .ZN(n381) );
  INV_X1 U430 ( .A(KEYINPUT105), .ZN(n382) );
  XOR2_X1 U431 ( .A(G116), .B(G107), .Z(n485) );
  INV_X1 U432 ( .A(G104), .ZN(n439) );
  XOR2_X1 U433 ( .A(G101), .B(G107), .Z(n418) );
  OR2_X1 U434 ( .A1(n673), .A2(n411), .ZN(n409) );
  NOR2_X1 U435 ( .A1(n697), .A2(n679), .ZN(n516) );
  BUF_X1 U436 ( .A(n680), .Z(n369) );
  OR2_X1 U437 ( .A1(n614), .A2(G902), .ZN(n482) );
  NOR2_X1 U438 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U439 ( .A(n414), .B(KEYINPUT77), .ZN(n413) );
  AND2_X1 U440 ( .A1(G953), .A2(G902), .ZN(n504) );
  XNOR2_X1 U441 ( .A(n699), .B(KEYINPUT80), .ZN(n580) );
  NOR2_X1 U442 ( .A1(n389), .A2(KEYINPUT106), .ZN(n386) );
  NAND2_X1 U443 ( .A1(n357), .A2(n370), .ZN(n387) );
  OR2_X1 U444 ( .A1(G237), .A2(G902), .ZN(n497) );
  XNOR2_X1 U445 ( .A(G116), .B(G137), .ZN(n473) );
  AND2_X1 U446 ( .A1(n597), .A2(n375), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n353), .B(G143), .ZN(n419) );
  XNOR2_X1 U448 ( .A(n489), .B(n488), .ZN(n402) );
  XNOR2_X1 U449 ( .A(n494), .B(n491), .ZN(n403) );
  XOR2_X1 U450 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n492) );
  NOR2_X1 U451 ( .A1(n525), .A2(KEYINPUT34), .ZN(n411) );
  XNOR2_X1 U452 ( .A(n523), .B(n522), .ZN(n673) );
  XNOR2_X1 U453 ( .A(n405), .B(KEYINPUT75), .ZN(n575) );
  NAND2_X1 U454 ( .A1(n406), .A2(n567), .ZN(n405) );
  INV_X1 U455 ( .A(G902), .ZN(n447) );
  XNOR2_X1 U456 ( .A(G128), .B(G119), .ZN(n452) );
  XNOR2_X1 U457 ( .A(KEYINPUT65), .B(n610), .ZN(n611) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n490), .B(n492), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n401) );
  AND2_X1 U461 ( .A1(n361), .A2(n663), .ZN(n587) );
  AND2_X1 U462 ( .A1(n521), .A2(n483), .ZN(n689) );
  NAND2_X1 U463 ( .A1(n559), .A2(n695), .ZN(n384) );
  BUF_X1 U464 ( .A(n517), .Z(n511) );
  XNOR2_X1 U465 ( .A(n614), .B(KEYINPUT62), .ZN(n615) );
  XNOR2_X1 U466 ( .A(n436), .B(n380), .ZN(n720) );
  XNOR2_X1 U467 ( .A(n445), .B(n381), .ZN(n380) );
  XNOR2_X1 U468 ( .A(n642), .B(n641), .ZN(n643) );
  BUF_X1 U469 ( .A(n638), .Z(n719) );
  XNOR2_X1 U470 ( .A(n479), .B(n446), .ZN(n714) );
  XNOR2_X1 U471 ( .A(n443), .B(n442), .ZN(n446) );
  XNOR2_X1 U472 ( .A(n490), .B(n418), .ZN(n443) );
  INV_X1 U473 ( .A(KEYINPUT35), .ZN(n371) );
  NAND2_X1 U474 ( .A1(n407), .A2(n359), .ZN(n372) );
  INV_X1 U475 ( .A(KEYINPUT32), .ZN(n539) );
  INV_X1 U476 ( .A(KEYINPUT107), .ZN(n397) );
  NOR2_X1 U477 ( .A1(n712), .A2(n711), .ZN(n713) );
  AND2_X1 U478 ( .A1(G210), .A2(n497), .ZN(n356) );
  AND2_X1 U479 ( .A1(n389), .A2(KEYINPUT106), .ZN(n357) );
  AND2_X1 U480 ( .A1(n394), .A2(n364), .ZN(n358) );
  AND2_X1 U481 ( .A1(n410), .A2(n417), .ZN(n359) );
  XOR2_X1 U482 ( .A(n560), .B(KEYINPUT38), .Z(n360) );
  AND2_X1 U483 ( .A1(n586), .A2(n695), .ZN(n361) );
  AND2_X1 U484 ( .A1(n684), .A2(n369), .ZN(n362) );
  AND2_X1 U485 ( .A1(n574), .A2(n360), .ZN(n363) );
  AND2_X1 U486 ( .A1(n534), .A2(n388), .ZN(n364) );
  XOR2_X1 U487 ( .A(KEYINPUT0), .B(KEYINPUT66), .Z(n365) );
  INV_X1 U488 ( .A(KEYINPUT106), .ZN(n388) );
  INV_X1 U489 ( .A(KEYINPUT34), .ZN(n412) );
  XNOR2_X1 U490 ( .A(KEYINPUT2), .B(KEYINPUT79), .ZN(n366) );
  XNOR2_X1 U491 ( .A(n367), .B(n455), .ZN(n460) );
  XNOR2_X1 U492 ( .A(n454), .B(n453), .ZN(n367) );
  NAND2_X1 U493 ( .A1(n368), .A2(n374), .ZN(n373) );
  XNOR2_X1 U494 ( .A(n377), .B(n573), .ZN(n368) );
  NAND2_X1 U495 ( .A1(n575), .A2(n363), .ZN(n562) );
  INV_X1 U496 ( .A(n662), .ZN(n392) );
  XNOR2_X1 U497 ( .A(n395), .B(KEYINPUT85), .ZN(n394) );
  INV_X1 U498 ( .A(n658), .ZN(n376) );
  INV_X1 U499 ( .A(n634), .ZN(n379) );
  INV_X1 U500 ( .A(n699), .ZN(n593) );
  XNOR2_X2 U501 ( .A(n496), .B(n356), .ZN(n559) );
  INV_X1 U502 ( .A(n653), .ZN(n393) );
  NAND2_X1 U503 ( .A1(n387), .A2(n385), .ZN(n530) );
  NOR2_X1 U504 ( .A1(n386), .A2(n358), .ZN(n385) );
  NAND2_X1 U505 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U506 ( .A1(n533), .A2(n589), .ZN(n395) );
  NAND2_X1 U507 ( .A1(n521), .A2(n535), .ZN(n523) );
  NAND2_X1 U508 ( .A1(n547), .A2(n396), .ZN(n548) );
  AND2_X1 U509 ( .A1(n546), .A2(n545), .ZN(n396) );
  XNOR2_X1 U510 ( .A(n533), .B(n397), .ZN(n398) );
  NAND2_X1 U511 ( .A1(n631), .A2(n751), .ZN(n543) );
  NOR2_X1 U512 ( .A1(n671), .A2(n495), .ZN(n612) );
  INV_X1 U513 ( .A(n555), .ZN(n406) );
  NAND2_X1 U514 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U515 ( .A1(n673), .A2(n412), .ZN(n408) );
  NAND2_X1 U516 ( .A1(n525), .A2(KEYINPUT34), .ZN(n410) );
  NOR2_X1 U517 ( .A1(n672), .A2(n413), .ZN(n675) );
  NAND2_X1 U518 ( .A1(n671), .A2(n366), .ZN(n414) );
  NOR2_X1 U519 ( .A1(n527), .A2(n526), .ZN(n417) );
  AND2_X1 U520 ( .A1(n668), .A2(n595), .ZN(n596) );
  INV_X1 U521 ( .A(KEYINPUT86), .ZN(n531) );
  NAND2_X1 U522 ( .A1(n724), .A2(n741), .ZN(n671) );
  XNOR2_X1 U523 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U524 ( .A(n736), .B(n441), .ZN(n442) );
  INV_X1 U525 ( .A(KEYINPUT63), .ZN(n619) );
  XNOR2_X1 U526 ( .A(n540), .B(n539), .ZN(n751) );
  XNOR2_X1 U527 ( .A(n419), .B(n486), .ZN(n423) );
  XOR2_X1 U528 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n421) );
  XNOR2_X1 U529 ( .A(G131), .B(G140), .ZN(n420) );
  XNOR2_X1 U530 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U531 ( .A(n423), .B(n422), .Z(n426) );
  XNOR2_X1 U532 ( .A(n493), .B(KEYINPUT10), .ZN(n737) );
  NOR2_X1 U533 ( .A1(G953), .A2(G237), .ZN(n472) );
  AND2_X1 U534 ( .A1(n472), .A2(G214), .ZN(n424) );
  XNOR2_X1 U535 ( .A(n737), .B(n424), .ZN(n425) );
  XNOR2_X1 U536 ( .A(n426), .B(n425), .ZN(n642) );
  NAND2_X1 U537 ( .A1(n642), .A2(n447), .ZN(n429) );
  XOR2_X1 U538 ( .A(G475), .B(KEYINPUT103), .Z(n427) );
  XNOR2_X1 U539 ( .A(KEYINPUT13), .B(n427), .ZN(n428) );
  XNOR2_X1 U540 ( .A(n429), .B(n428), .ZN(n527) );
  XOR2_X1 U541 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n431) );
  XNOR2_X1 U542 ( .A(G122), .B(KEYINPUT9), .ZN(n430) );
  XNOR2_X1 U543 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X2 U544 ( .A(G143), .B(G128), .ZN(n489) );
  NAND2_X1 U545 ( .A1(n742), .A2(G234), .ZN(n433) );
  XNOR2_X1 U546 ( .A(n434), .B(n433), .ZN(n449) );
  NAND2_X1 U547 ( .A1(n449), .A2(G217), .ZN(n435) );
  XNOR2_X1 U548 ( .A(n485), .B(n435), .ZN(n436) );
  NOR2_X1 U549 ( .A1(G902), .A2(n720), .ZN(n437) );
  XNOR2_X1 U550 ( .A(n437), .B(G478), .ZN(n526) );
  INV_X1 U551 ( .A(n526), .ZN(n438) );
  AND2_X1 U552 ( .A1(n527), .A2(n438), .ZN(n665) );
  NOR2_X1 U553 ( .A1(n663), .A2(n665), .ZN(n699) );
  XOR2_X1 U554 ( .A(KEYINPUT68), .B(G110), .Z(n490) );
  XNOR2_X1 U555 ( .A(n457), .B(KEYINPUT95), .ZN(n736) );
  NAND2_X1 U556 ( .A1(G227), .A2(n742), .ZN(n440) );
  XNOR2_X1 U557 ( .A(KEYINPUT4), .B(G131), .ZN(n444) );
  NAND2_X1 U558 ( .A1(n714), .A2(n447), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n570), .B(KEYINPUT1), .ZN(n519) );
  NAND2_X1 U560 ( .A1(n449), .A2(G221), .ZN(n455) );
  XNOR2_X1 U561 ( .A(G110), .B(KEYINPUT23), .ZN(n451) );
  XNOR2_X1 U562 ( .A(KEYINPUT24), .B(KEYINPUT97), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n451), .B(n450), .ZN(n454) );
  XNOR2_X1 U564 ( .A(n452), .B(KEYINPUT98), .ZN(n453) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(KEYINPUT96), .ZN(n456) );
  XNOR2_X1 U566 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n737), .B(n458), .ZN(n459) );
  XNOR2_X1 U568 ( .A(n460), .B(n459), .ZN(n636) );
  XOR2_X1 U569 ( .A(n461), .B(KEYINPUT89), .Z(n495) );
  NAND2_X1 U570 ( .A1(n495), .A2(G234), .ZN(n462) );
  XNOR2_X1 U571 ( .A(n462), .B(KEYINPUT20), .ZN(n466) );
  NAND2_X1 U572 ( .A1(n466), .A2(G217), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n463), .B(KEYINPUT25), .ZN(n464) );
  NAND2_X1 U574 ( .A1(n466), .A2(G221), .ZN(n469) );
  INV_X1 U575 ( .A(KEYINPUT99), .ZN(n467) );
  XNOR2_X1 U576 ( .A(n467), .B(KEYINPUT21), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n469), .B(n468), .ZN(n679) );
  NOR2_X2 U578 ( .A1(n680), .A2(n679), .ZN(n677) );
  NAND2_X1 U579 ( .A1(n519), .A2(n677), .ZN(n470) );
  NAND2_X1 U580 ( .A1(n472), .A2(G210), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U582 ( .A(KEYINPUT101), .B(KEYINPUT5), .ZN(n475) );
  XNOR2_X1 U583 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U584 ( .A(n484), .B(n477), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n479), .B(n478), .ZN(n614) );
  INV_X1 U586 ( .A(KEYINPUT70), .ZN(n480) );
  XNOR2_X1 U587 ( .A(n480), .B(G472), .ZN(n481) );
  XNOR2_X2 U588 ( .A(n482), .B(n481), .ZN(n684) );
  INV_X1 U589 ( .A(n684), .ZN(n483) );
  NAND2_X1 U590 ( .A1(G224), .A2(n742), .ZN(n488) );
  XNOR2_X1 U591 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n491) );
  INV_X1 U592 ( .A(n493), .ZN(n494) );
  INV_X1 U593 ( .A(n495), .ZN(n609) );
  NAND2_X1 U594 ( .A1(n624), .A2(n495), .ZN(n496) );
  NAND2_X1 U595 ( .A1(G214), .A2(n497), .ZN(n499) );
  INV_X1 U596 ( .A(KEYINPUT91), .ZN(n498) );
  INV_X1 U597 ( .A(KEYINPUT19), .ZN(n500) );
  NAND2_X1 U598 ( .A1(G234), .A2(G237), .ZN(n501) );
  XNOR2_X1 U599 ( .A(n501), .B(KEYINPUT92), .ZN(n502) );
  XNOR2_X1 U600 ( .A(KEYINPUT14), .B(n502), .ZN(n505) );
  NAND2_X1 U601 ( .A1(G952), .A2(n505), .ZN(n710) );
  NOR2_X1 U602 ( .A1(G953), .A2(n710), .ZN(n503) );
  XOR2_X1 U603 ( .A(KEYINPUT93), .B(n503), .Z(n552) );
  NAND2_X1 U604 ( .A1(n505), .A2(n504), .ZN(n549) );
  NOR2_X1 U605 ( .A1(G898), .A2(n549), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n506), .B(KEYINPUT94), .ZN(n507) );
  NAND2_X1 U607 ( .A1(n689), .A2(n511), .ZN(n510) );
  XNOR2_X1 U608 ( .A(n510), .B(KEYINPUT31), .ZN(n662) );
  NAND2_X1 U609 ( .A1(n511), .A2(n684), .ZN(n513) );
  NAND2_X1 U610 ( .A1(n677), .A2(n570), .ZN(n512) );
  XNOR2_X1 U611 ( .A(n512), .B(KEYINPUT100), .ZN(n555) );
  INV_X1 U612 ( .A(KEYINPUT6), .ZN(n515) );
  NAND2_X1 U613 ( .A1(n526), .A2(n527), .ZN(n697) );
  NOR2_X2 U614 ( .A1(n538), .A2(n520), .ZN(n533) );
  INV_X1 U615 ( .A(n369), .ZN(n534) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n528) );
  INV_X1 U617 ( .A(n589), .ZN(n535) );
  INV_X1 U618 ( .A(KEYINPUT33), .ZN(n522) );
  BUF_X1 U619 ( .A(n524), .Z(n525) );
  NAND2_X1 U620 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U621 ( .A(n532), .B(n531), .ZN(n547) );
  NOR2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n520), .A2(n536), .ZN(n537) );
  NOR2_X1 U624 ( .A1(n538), .A2(n537), .ZN(n540) );
  NOR2_X1 U625 ( .A1(n543), .A2(KEYINPUT44), .ZN(n541) );
  XNOR2_X1 U626 ( .A(n542), .B(KEYINPUT69), .ZN(n546) );
  BUF_X1 U627 ( .A(n543), .Z(n544) );
  NAND2_X1 U628 ( .A1(n544), .A2(KEYINPUT44), .ZN(n545) );
  XNOR2_X2 U629 ( .A(n548), .B(KEYINPUT45), .ZN(n724) );
  XNOR2_X1 U630 ( .A(KEYINPUT108), .B(n549), .ZN(n550) );
  NOR2_X1 U631 ( .A1(G900), .A2(n550), .ZN(n551) );
  NOR2_X1 U632 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U633 ( .A(KEYINPUT76), .ZN(n553) );
  XNOR2_X1 U634 ( .A(n554), .B(n553), .ZN(n567) );
  INV_X1 U635 ( .A(n695), .ZN(n556) );
  OR2_X1 U636 ( .A1(n684), .A2(n556), .ZN(n558) );
  XNOR2_X1 U637 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n557) );
  XNOR2_X1 U638 ( .A(n558), .B(n557), .ZN(n574) );
  BUF_X1 U639 ( .A(n559), .Z(n560) );
  XNOR2_X1 U640 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n561) );
  NAND2_X1 U641 ( .A1(n599), .A2(n663), .ZN(n564) );
  INV_X1 U642 ( .A(KEYINPUT40), .ZN(n563) );
  XNOR2_X1 U643 ( .A(n564), .B(n563), .ZN(n634) );
  NAND2_X1 U644 ( .A1(n360), .A2(n695), .ZN(n700) );
  NOR2_X1 U645 ( .A1(n700), .A2(n697), .ZN(n565) );
  XNOR2_X1 U646 ( .A(KEYINPUT41), .B(n565), .ZN(n693) );
  INV_X1 U647 ( .A(n679), .ZN(n566) );
  AND2_X1 U648 ( .A1(n567), .A2(n566), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n586), .A2(n369), .ZN(n568) );
  NOR2_X1 U650 ( .A1(n568), .A2(n684), .ZN(n569) );
  XNOR2_X1 U651 ( .A(n569), .B(KEYINPUT28), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n571), .A2(n570), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n693), .A2(n582), .ZN(n572) );
  XNOR2_X1 U654 ( .A(n572), .B(KEYINPUT42), .ZN(n752) );
  INV_X1 U655 ( .A(KEYINPUT46), .ZN(n573) );
  AND2_X1 U656 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n576), .A2(n560), .ZN(n578) );
  INV_X1 U658 ( .A(KEYINPUT110), .ZN(n577) );
  XNOR2_X1 U659 ( .A(n578), .B(n577), .ZN(n579) );
  AND2_X1 U660 ( .A1(n579), .A2(n417), .ZN(n658) );
  NOR2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n659) );
  NAND2_X1 U662 ( .A1(n583), .A2(n659), .ZN(n585) );
  INV_X1 U663 ( .A(KEYINPUT71), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n585), .B(n584), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n587), .A2(n369), .ZN(n588) );
  OR2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n600) );
  INV_X1 U667 ( .A(n560), .ZN(n602) );
  OR2_X1 U668 ( .A1(n600), .A2(n602), .ZN(n591) );
  INV_X1 U669 ( .A(KEYINPUT36), .ZN(n590) );
  XNOR2_X1 U670 ( .A(n591), .B(n590), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n520), .A2(n592), .ZN(n668) );
  NAND2_X1 U672 ( .A1(n659), .A2(n593), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n594), .A2(KEYINPUT47), .ZN(n595) );
  XNOR2_X1 U674 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n665), .ZN(n632) );
  OR2_X1 U676 ( .A1(n520), .A2(n600), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT43), .ZN(n603) );
  AND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n669) );
  INV_X1 U679 ( .A(n669), .ZN(n604) );
  AND2_X1 U680 ( .A1(n632), .A2(n604), .ZN(n605) );
  AND2_X1 U681 ( .A1(n741), .A2(KEYINPUT2), .ZN(n607) );
  XNOR2_X2 U682 ( .A(n608), .B(KEYINPUT74), .ZN(n672) );
  NAND2_X1 U683 ( .A1(n609), .A2(KEYINPUT2), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X4 U685 ( .A1(n672), .A2(n613), .ZN(n638) );
  NAND2_X1 U686 ( .A1(n638), .A2(G472), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n618) );
  INV_X1 U688 ( .A(G952), .ZN(n617) );
  AND2_X1 U689 ( .A1(n617), .A2(G953), .ZN(n723) );
  NOR2_X2 U690 ( .A1(n618), .A2(n723), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(G57) );
  NAND2_X1 U692 ( .A1(n638), .A2(G210), .ZN(n626) );
  XOR2_X1 U693 ( .A(KEYINPUT87), .B(KEYINPUT78), .Z(n622) );
  XNOR2_X1 U694 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U698 ( .A1(n627), .A2(n723), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(KEYINPUT122), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT56), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(G51) );
  XNOR2_X1 U702 ( .A(n631), .B(G110), .ZN(G12) );
  XNOR2_X1 U703 ( .A(n632), .B(G134), .ZN(G36) );
  XOR2_X1 U704 ( .A(n633), .B(G101), .Z(G3) );
  XOR2_X1 U705 ( .A(n634), .B(G131), .Z(G33) );
  NAND2_X1 U706 ( .A1(n719), .A2(G217), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X1 U708 ( .A1(n637), .A2(n723), .ZN(G66) );
  NAND2_X1 U709 ( .A1(n638), .A2(G475), .ZN(n644) );
  XOR2_X1 U710 ( .A(KEYINPUT88), .B(KEYINPUT123), .Z(n640) );
  XNOR2_X1 U711 ( .A(KEYINPUT59), .B(KEYINPUT64), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U714 ( .A1(n645), .A2(n723), .ZN(n647) );
  XNOR2_X1 U715 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G60) );
  XOR2_X1 U717 ( .A(G104), .B(KEYINPUT111), .Z(n649) );
  NAND2_X1 U718 ( .A1(n663), .A2(n354), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n651) );
  XNOR2_X1 U721 ( .A(G107), .B(KEYINPUT26), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(n652), .Z(n655) );
  NAND2_X1 U724 ( .A1(n665), .A2(n354), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(G9) );
  XOR2_X1 U726 ( .A(G128), .B(KEYINPUT29), .Z(n657) );
  NAND2_X1 U727 ( .A1(n665), .A2(n659), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(G30) );
  XOR2_X1 U729 ( .A(G143), .B(n658), .Z(G45) );
  NAND2_X1 U730 ( .A1(n659), .A2(n663), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(KEYINPUT114), .ZN(n661) );
  XNOR2_X1 U732 ( .A(G146), .B(n661), .ZN(G48) );
  NAND2_X1 U733 ( .A1(n662), .A2(n663), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(n353), .ZN(G15) );
  NAND2_X1 U735 ( .A1(n662), .A2(n665), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(G116), .ZN(G18) );
  XOR2_X1 U737 ( .A(G125), .B(KEYINPUT37), .Z(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G27) );
  XNOR2_X1 U739 ( .A(G140), .B(n669), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n670), .B(KEYINPUT115), .ZN(G42) );
  BUF_X1 U741 ( .A(n673), .Z(n703) );
  NOR2_X1 U742 ( .A1(n703), .A2(n693), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n676), .A2(n742), .ZN(n712) );
  NOR2_X1 U744 ( .A1(n520), .A2(n677), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT50), .ZN(n687) );
  NAND2_X1 U746 ( .A1(n369), .A2(n679), .ZN(n683) );
  XNOR2_X1 U747 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(KEYINPUT116), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n688), .B(KEYINPUT118), .ZN(n690) );
  NOR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U754 ( .A(KEYINPUT51), .B(n691), .Z(n692) );
  NOR2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U756 ( .A(KEYINPUT119), .B(n694), .Z(n706) );
  NOR2_X1 U757 ( .A1(n360), .A2(n695), .ZN(n696) );
  NOR2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U759 ( .A(n698), .B(KEYINPUT120), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U764 ( .A(n707), .B(KEYINPUT121), .Z(n708) );
  XNOR2_X1 U765 ( .A(KEYINPUT52), .B(n708), .ZN(n709) );
  NOR2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U768 ( .A1(n719), .A2(G469), .ZN(n717) );
  XOR2_X1 U769 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XOR2_X1 U770 ( .A(n715), .B(n714), .Z(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n723), .A2(n718), .ZN(G54) );
  NAND2_X1 U773 ( .A1(n719), .A2(G478), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n723), .A2(n722), .ZN(G63) );
  BUF_X1 U776 ( .A(n724), .Z(n725) );
  NAND2_X1 U777 ( .A1(n742), .A2(n725), .ZN(n729) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n726) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n726), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n727), .A2(G898), .ZN(n728) );
  NAND2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n730), .B(G110), .ZN(n732) );
  NOR2_X1 U783 ( .A1(n742), .A2(G898), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n735) );
  XOR2_X1 U786 ( .A(KEYINPUT125), .B(n735), .Z(G69) );
  XNOR2_X1 U787 ( .A(n736), .B(KEYINPUT126), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n739) );
  XOR2_X1 U789 ( .A(n740), .B(n739), .Z(n744) );
  XNOR2_X1 U790 ( .A(n741), .B(n744), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n748) );
  XOR2_X1 U792 ( .A(G227), .B(n744), .Z(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G953), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U796 ( .A(n749), .B(G122), .Z(n750) );
  XNOR2_X1 U797 ( .A(n750), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U798 ( .A(G119), .B(n751), .ZN(G21) );
  XOR2_X1 U799 ( .A(G137), .B(n752), .Z(G39) );
endmodule

