//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n466), .A2(new_n463), .A3(G101), .A4(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n463), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n470), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n463), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n485), .B1(new_n488), .B2(G136), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT69), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n463), .C1(new_n469), .C2(new_n470), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n486), .A2(new_n499), .A3(G138), .A4(new_n463), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(new_n502), .A3(KEYINPUT5), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n511), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT7), .Z(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(G51), .B2(new_n514), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n508), .A2(new_n516), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n510), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n514), .A2(G52), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT71), .B(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n517), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n505), .A2(new_n507), .ZN(new_n537));
  INV_X1    g112(.A(new_n503), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n535), .B(new_n536), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n510), .B1(new_n542), .B2(KEYINPUT72), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n508), .A2(G81), .A3(new_n516), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n514), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT73), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n541), .A2(new_n543), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT75), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  AND2_X1   g133(.A1(KEYINPUT6), .A2(G651), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT6), .A2(G651), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n516), .A2(G53), .A3(G543), .A4(new_n562), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n539), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n524), .B2(G91), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n558), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n562), .B1(new_n514), .B2(G53), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n561), .A2(new_n563), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT77), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n508), .A2(G91), .A3(new_n516), .ZN(new_n580));
  INV_X1    g155(.A(new_n570), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n508), .B2(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n582), .B2(new_n510), .ZN(new_n583));
  NOR3_X1   g158(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n574), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G166), .ZN(G303));
  OAI21_X1  g162(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n508), .A2(G87), .A3(new_n516), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n514), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n514), .A2(G48), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n510), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n537), .A2(G86), .A3(new_n538), .A4(new_n516), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n508), .A2(KEYINPUT79), .A3(G86), .A4(new_n516), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n510), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n514), .A2(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n517), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n603), .B2(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n508), .A2(G92), .A3(new_n516), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT10), .Z(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT81), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n539), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT82), .Z(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G299), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n626), .ZN(G297));
  XNOR2_X1  g202(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n620), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n543), .A2(new_n541), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n547), .A2(new_n549), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n625), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n619), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n479), .A2(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n463), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n638), .B1(new_n639), .B2(new_n640), .C1(new_n641), .C2(new_n487), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT84), .Z(G156));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n656), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n671), .B1(new_n672), .B2(new_n669), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI22_X1  g251(.A1(new_n670), .A2(new_n672), .B1(new_n676), .B2(KEYINPUT87), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(KEYINPUT87), .B2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(new_n671), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n672), .A3(new_n669), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n674), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n688), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  MUX2_X1   g269(.A(new_n688), .B(new_n693), .S(new_n694), .Z(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n688), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n699), .B1(new_n695), .B2(new_n698), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n686), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(new_n686), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(new_n705), .A3(new_n700), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n703), .B2(new_n706), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(G166), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G22), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(G6), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n600), .B2(new_n711), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n713), .A2(new_n714), .ZN(new_n720));
  MUX2_X1   g295(.A(G23), .B(G288), .S(G16), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NOR4_X1   g298(.A1(new_n715), .A2(new_n719), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n711), .A2(G24), .ZN(new_n728));
  INV_X1    g303(.A(G290), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n711), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G1986), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G1986), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n479), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n463), .A2(G107), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(G131), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n733), .B1(new_n734), .B2(new_n735), .C1(new_n736), .C2(new_n487), .ZN(new_n737));
  MUX2_X1   g312(.A(G25), .B(new_n737), .S(G29), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT35), .B(G1991), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n731), .A2(new_n732), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n726), .A2(new_n727), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G32), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n479), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G141), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n487), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n759), .B2(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT24), .B2(new_n759), .ZN(new_n761));
  INV_X1    g336(.A(G160), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n746), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT96), .Z(new_n766));
  XOR2_X1   g341(.A(KEYINPUT31), .B(G11), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT30), .B(G28), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n767), .B1(new_n746), .B2(new_n768), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n769), .B1(new_n746), .B2(new_n642), .C1(new_n763), .C2(new_n764), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G21), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G168), .B2(G16), .ZN(new_n772));
  NOR2_X1   g347(.A1(G27), .A2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(G29), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n772), .A2(G1966), .B1(G2078), .B2(new_n774), .ZN(new_n775));
  OR4_X1    g350(.A1(new_n758), .A2(new_n766), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n711), .A2(G5), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G171), .B2(new_n711), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1961), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n746), .A2(G26), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT28), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n488), .A2(G140), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n479), .A2(G128), .ZN(new_n783));
  OR2_X1    g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n781), .B1(new_n787), .B2(new_n746), .ZN(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n772), .A2(G1966), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n774), .A2(G2078), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n550), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1341), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n776), .A2(new_n779), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G29), .A2(G35), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G162), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT29), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G2090), .ZN(new_n801));
  NOR2_X1   g376(.A1(G29), .A2(G33), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  INV_X1    g378(.A(G127), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n477), .B2(new_n478), .ZN(new_n805));
  AND2_X1   g380(.A1(G115), .A2(G2104), .ZN(new_n806));
  OAI21_X1  g381(.A(G2105), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n811));
  NAND2_X1  g386(.A1(G103), .A2(G2104), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G2105), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n488), .A2(G139), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n803), .B1(new_n816), .B2(new_n746), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G2072), .Z(new_n818));
  NOR2_X1   g393(.A1(G4), .A2(G16), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n620), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT93), .B(G1348), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  AOI211_X1 g397(.A(new_n818), .B(new_n822), .C1(new_n800), .C2(G2090), .ZN(new_n823));
  NAND2_X1  g398(.A1(G299), .A2(G16), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n711), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT23), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G1956), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n797), .A2(new_n801), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n745), .A2(new_n830), .ZN(G311));
  INV_X1    g406(.A(G311), .ZN(G150));
  AND2_X1   g407(.A1(G80), .A2(G543), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n508), .B2(G67), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n835));
  OAI21_X1  g410(.A(G651), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n537), .A2(G67), .A3(new_n538), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n837), .A2(KEYINPUT98), .A3(new_n833), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT99), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT98), .B1(new_n837), .B2(new_n833), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n834), .A2(new_n835), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(G651), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n514), .A2(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n517), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n839), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n620), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n848), .A2(new_n633), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n840), .A2(new_n841), .A3(G651), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n846), .B1(new_n855), .B2(KEYINPUT99), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n550), .A3(new_n843), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  INV_X1    g435(.A(G860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n859), .B2(KEYINPUT39), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n850), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT100), .ZN(G145));
  NAND2_X1  g439(.A1(new_n479), .A2(G130), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n463), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G142), .B2(new_n488), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n645), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n737), .ZN(new_n871));
  INV_X1    g446(.A(new_n755), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n816), .A2(new_n872), .A3(KEYINPUT101), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n816), .B2(KEYINPUT101), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n787), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n755), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n786), .A3(new_n873), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(G164), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G164), .B1(new_n876), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n879), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n498), .A2(new_n500), .ZN(new_n885));
  INV_X1    g460(.A(new_n496), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n870), .B(new_n737), .Z(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n880), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G162), .B(new_n642), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G160), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n892), .B(new_n762), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n888), .A2(new_n889), .A3(new_n880), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .A4(new_n883), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT103), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(G395));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT104), .B1(new_n574), .B2(new_n584), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT78), .B1(new_n579), .B2(new_n583), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n569), .A2(new_n573), .A3(new_n558), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n619), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n620), .B(KEYINPUT104), .C1(new_n574), .C2(new_n584), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n848), .A2(new_n633), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n550), .B1(new_n856), .B2(new_n843), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n635), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n854), .B(new_n857), .C1(G559), .C2(new_n619), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n913), .A2(new_n914), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(KEYINPUT105), .A3(new_n920), .A4(new_n921), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n922), .B2(new_n915), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n917), .A2(KEYINPUT106), .A3(new_n922), .A4(new_n923), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n907), .A2(new_n926), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(new_n931), .A3(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT107), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n729), .A2(G305), .ZN(new_n936));
  NOR2_X1   g511(.A1(G290), .A2(new_n600), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(G166), .B(G288), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n936), .B2(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT42), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n933), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n944), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n946), .A2(new_n934), .A3(KEYINPUT107), .ZN(new_n947));
  OAI21_X1  g522(.A(G868), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n848), .A2(new_n625), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(G295));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n949), .ZN(G331));
  XOR2_X1   g526(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(G301), .A2(G168), .ZN(new_n954));
  NAND2_X1  g529(.A1(G171), .A2(G286), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n918), .B2(new_n919), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n854), .A2(new_n857), .A3(new_n955), .A4(new_n954), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n959), .B2(new_n915), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n917), .A3(new_n923), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n958), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n927), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n961), .A3(new_n964), .A4(new_n943), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n968));
  INV_X1    g543(.A(new_n943), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n953), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n959), .A2(new_n917), .A3(new_n923), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n959), .A2(new_n915), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(new_n966), .A3(new_n965), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n952), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n967), .A2(new_n953), .A3(new_n970), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT44), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n887), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n472), .A2(new_n475), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n987), .A2(new_n988), .A3(new_n755), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT112), .ZN(new_n990));
  INV_X1    g565(.A(new_n987), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n786), .B(G2067), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n987), .A2(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT111), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(new_n872), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n737), .A2(new_n740), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n737), .A2(new_n740), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OR3_X1    g575(.A1(G290), .A2(G1986), .A3(new_n987), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT48), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n995), .B(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n991), .B1(new_n992), .B2(new_n872), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1005), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n787), .A2(new_n789), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n993), .A2(new_n996), .ZN(new_n1011));
  INV_X1    g586(.A(new_n999), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(new_n991), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT126), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1008), .A2(new_n1007), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT126), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n991), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1003), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n887), .A2(new_n1022), .A3(new_n982), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1023), .A3(new_n986), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n885), .B2(new_n886), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n986), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1024), .A2(new_n821), .B1(new_n1027), .B2(new_n789), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n619), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n828), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n984), .B1(G164), .B2(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n986), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n579), .A2(new_n1036), .A3(new_n583), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n583), .A2(KEYINPUT120), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n564), .A2(new_n565), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n580), .C1(new_n582), .C2(new_n510), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1029), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G160), .A2(G40), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1956), .B1(new_n1046), .B2(new_n1023), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1034), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT121), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1030), .A2(new_n1050), .A3(new_n1034), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1051), .A3(new_n1043), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1031), .A2(new_n1032), .A3(new_n986), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1055), .A2(new_n1033), .B1(new_n1024), .B2(new_n828), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1042), .A2(new_n1036), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1037), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1052), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1054), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n986), .B1(new_n1025), .B2(new_n1022), .ZN(new_n1065));
  NOR3_X1   g640(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n821), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1027), .A2(new_n789), .ZN(new_n1068));
  AND4_X1   g643(.A1(KEYINPUT60), .A2(new_n1067), .A3(new_n619), .A4(new_n1068), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1028), .A2(KEYINPUT60), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n619), .B1(new_n1028), .B2(KEYINPUT60), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1061), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1031), .A2(new_n1032), .A3(new_n988), .A4(new_n986), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  AOI22_X1  g650(.A1(new_n1074), .A2(KEYINPUT122), .B1(new_n1026), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1055), .A2(new_n1077), .A3(new_n988), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n633), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT59), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1053), .B1(new_n1073), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1031), .A2(new_n1032), .A3(new_n986), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(G2078), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1045), .B1(new_n983), .B2(new_n984), .ZN(new_n1085));
  INV_X1    g660(.A(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(KEYINPUT53), .A3(new_n1086), .A4(new_n1032), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1024), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1084), .A2(new_n1087), .A3(G301), .A4(new_n1089), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(KEYINPUT54), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT124), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  AND4_X1   g670(.A1(new_n1086), .A2(new_n1031), .A3(new_n1032), .A4(new_n986), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(KEYINPUT53), .B1(new_n1088), .B2(new_n1024), .ZN(new_n1097));
  AOI21_X1  g672(.A(G301), .B1(new_n1097), .B2(new_n1084), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1092), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G286), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n1101), .B2(KEYINPUT123), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT117), .B(G2084), .Z(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1104), .A2(new_n1105), .B1(new_n1083), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1101), .B(new_n1103), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1105), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1055), .A2(G1966), .B1(new_n1024), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(G8), .B(new_n1102), .C1(new_n1111), .C2(G286), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(G8), .A3(G286), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n594), .A2(new_n599), .A3(G1981), .ZN(new_n1116));
  INV_X1    g691(.A(G1981), .ZN(new_n1117));
  INV_X1    g692(.A(new_n592), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n537), .A2(G61), .A3(new_n538), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G73), .A2(G543), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1121), .B2(G651), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(new_n595), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1115), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT49), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT49), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1115), .B(new_n1126), .C1(new_n1116), .C2(new_n1123), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1108), .B1(new_n1025), .B2(new_n986), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT113), .B(G1971), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1083), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G2090), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1021), .A2(new_n1023), .A3(new_n1132), .A4(new_n986), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT55), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(G166), .B2(new_n1108), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT55), .B(G8), .C1(new_n511), .C2(new_n519), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(G8), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1976), .ZN(new_n1140));
  OR2_X1    g715(.A1(G288), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT52), .B1(G288), .B2(new_n1140), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1128), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1128), .A2(new_n1141), .A3(KEYINPUT114), .A4(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1145), .A2(new_n1146), .B1(KEYINPUT52), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1129), .A2(new_n1139), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1108), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT116), .B1(new_n1150), .B2(new_n1138), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1138), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1104), .A2(new_n1132), .B1(new_n1083), .B2(new_n1130), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1152), .B(new_n1153), .C1(new_n1154), .C2(new_n1108), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1100), .A2(new_n1114), .A3(new_n1149), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1081), .A2(new_n1094), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(G288), .A2(G1976), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1116), .B1(new_n1129), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1128), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1129), .A2(new_n1148), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1160), .A2(new_n1161), .B1(new_n1162), .B2(new_n1139), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1107), .A2(new_n1108), .A3(G286), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1149), .A2(new_n1156), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(new_n1153), .A3(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1170), .A2(new_n1149), .A3(KEYINPUT63), .A4(new_n1164), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1163), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1114), .A2(KEYINPUT62), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1114), .A2(KEYINPUT62), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1098), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1158), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(G290), .A2(G1986), .A3(new_n991), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1001), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT110), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n997), .A2(new_n1000), .A3(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1177), .A2(KEYINPUT125), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT125), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1020), .B1(new_n1182), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g759(.A1(new_n971), .A2(new_n976), .ZN(new_n1186));
  NOR3_X1   g760(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1187));
  OAI21_X1  g761(.A(new_n1187), .B1(new_n708), .B2(new_n709), .ZN(new_n1188));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g764(.A(new_n1187), .B(KEYINPUT127), .C1(new_n708), .C2(new_n709), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n902), .B1(new_n894), .B2(new_n899), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1186), .A2(new_n1195), .ZN(G308));
  OAI221_X1 g770(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .C1(new_n971), .C2(new_n976), .ZN(G225));
endmodule


