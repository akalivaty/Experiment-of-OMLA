

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748;

  XNOR2_X1 U359 ( .A(n338), .B(n337), .ZN(n629) );
  INV_X1 U360 ( .A(KEYINPUT32), .ZN(n337) );
  AND2_X1 U361 ( .A1(n553), .A2(n552), .ZN(n663) );
  XNOR2_X1 U362 ( .A(n388), .B(n434), .ZN(n524) );
  XNOR2_X1 U363 ( .A(G116), .B(KEYINPUT3), .ZN(n407) );
  AND2_X1 U364 ( .A1(n378), .A2(n354), .ZN(n344) );
  NAND2_X2 U365 ( .A1(n372), .A2(n488), .ZN(n342) );
  XNOR2_X2 U366 ( .A(n364), .B(n484), .ZN(n372) );
  XNOR2_X2 U367 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X2 U368 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n362) );
  AND2_X2 U369 ( .A1(n610), .A2(n740), .ZN(n672) );
  XNOR2_X1 U370 ( .A(n560), .B(n559), .ZN(n610) );
  NAND2_X1 U371 ( .A1(n612), .A2(n676), .ZN(n345) );
  XNOR2_X2 U372 ( .A(n544), .B(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U373 ( .A1(n536), .A2(n375), .ZN(n338) );
  XNOR2_X2 U374 ( .A(n632), .B(n426), .ZN(n617) );
  XOR2_X2 U375 ( .A(n566), .B(KEYINPUT28), .Z(n568) );
  XOR2_X2 U376 ( .A(n634), .B(n633), .Z(n358) );
  BUF_X2 U377 ( .A(n370), .Z(n339) );
  XNOR2_X2 U378 ( .A(n400), .B(G143), .ZN(n388) );
  XNOR2_X2 U379 ( .A(n444), .B(G110), .ZN(n385) );
  NOR2_X1 U380 ( .A1(n672), .A2(KEYINPUT2), .ZN(n607) );
  NOR2_X2 U381 ( .A1(n586), .A2(n659), .ZN(n602) );
  XOR2_X2 U382 ( .A(KEYINPUT10), .B(n481), .Z(n501) );
  XNOR2_X1 U383 ( .A(G137), .B(G101), .ZN(n416) );
  XNOR2_X1 U384 ( .A(n524), .B(n397), .ZN(n735) );
  INV_X1 U385 ( .A(G953), .ZN(n741) );
  NOR2_X2 U386 ( .A1(n376), .A2(n347), .ZN(n402) );
  NOR2_X2 U387 ( .A1(n541), .A2(n540), .ZN(n543) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n436) );
  XNOR2_X1 U389 ( .A(n595), .B(KEYINPUT41), .ZN(n708) );
  AND2_X1 U390 ( .A1(n590), .A2(n346), .ZN(n669) );
  AND2_X1 U391 ( .A1(n707), .A2(KEYINPUT34), .ZN(n347) );
  NOR2_X1 U392 ( .A1(n391), .A2(n545), .ZN(n472) );
  XNOR2_X1 U393 ( .A(n517), .B(n516), .ZN(n553) );
  XNOR2_X1 U394 ( .A(n374), .B(n373), .ZN(n567) );
  XNOR2_X1 U395 ( .A(n514), .B(n513), .ZN(n634) );
  XNOR2_X1 U396 ( .A(n735), .B(G146), .ZN(n442) );
  XNOR2_X1 U397 ( .A(n398), .B(n480), .ZN(n397) );
  XNOR2_X1 U398 ( .A(n435), .B(KEYINPUT4), .ZN(n480) );
  XNOR2_X1 U399 ( .A(G107), .B(G104), .ZN(n443) );
  INV_X1 U400 ( .A(KEYINPUT66), .ZN(n435) );
  INV_X2 U401 ( .A(G125), .ZN(n455) );
  INV_X1 U402 ( .A(G128), .ZN(n400) );
  XNOR2_X2 U403 ( .A(n340), .B(n491), .ZN(n587) );
  NAND2_X2 U404 ( .A1(n341), .A2(n342), .ZN(n340) );
  AND2_X2 U405 ( .A1(n428), .A2(n348), .ZN(n341) );
  OR2_X2 U406 ( .A1(n638), .A2(n429), .ZN(n428) );
  NAND2_X1 U407 ( .A1(n355), .A2(n342), .ZN(n581) );
  XNOR2_X2 U408 ( .A(n587), .B(n356), .ZN(n569) );
  BUF_X1 U409 ( .A(n536), .Z(n343) );
  AND2_X1 U410 ( .A1(n378), .A2(n354), .ZN(n740) );
  NAND2_X1 U411 ( .A1(n612), .A2(n676), .ZN(n632) );
  AND2_X2 U412 ( .A1(n569), .A2(n567), .ZN(n421) );
  BUF_X1 U413 ( .A(n537), .Z(n346) );
  XNOR2_X1 U414 ( .A(n567), .B(KEYINPUT1), .ZN(n537) );
  NOR2_X2 U415 ( .A1(n690), .A2(n370), .ZN(n577) );
  XNOR2_X2 U416 ( .A(n475), .B(n473), .ZN(n379) );
  XNOR2_X2 U417 ( .A(n439), .B(n438), .ZN(n474) );
  XOR2_X1 U418 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n504) );
  XNOR2_X1 U419 ( .A(n399), .B(KEYINPUT67), .ZN(n502) );
  INV_X1 U420 ( .A(G131), .ZN(n399) );
  INV_X1 U421 ( .A(n485), .ZN(n431) );
  XNOR2_X1 U422 ( .A(KEYINPUT16), .B(G122), .ZN(n473) );
  INV_X1 U423 ( .A(G237), .ZN(n486) );
  NAND2_X1 U424 ( .A1(n619), .A2(n487), .ZN(n441) );
  INV_X1 U425 ( .A(G469), .ZN(n373) );
  XOR2_X1 U426 ( .A(KEYINPUT11), .B(G122), .Z(n512) );
  NOR2_X1 U427 ( .A1(n500), .A2(KEYINPUT34), .ZN(n404) );
  INV_X1 U428 ( .A(KEYINPUT22), .ZN(n424) );
  XNOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n477) );
  XNOR2_X1 U430 ( .A(n505), .B(n433), .ZN(n506) );
  XNOR2_X1 U431 ( .A(KEYINPUT97), .B(KEYINPUT12), .ZN(n503) );
  XNOR2_X1 U432 ( .A(G143), .B(G113), .ZN(n509) );
  NAND2_X1 U433 ( .A1(n679), .A2(n564), .ZN(n419) );
  NAND2_X1 U434 ( .A1(n485), .A2(n488), .ZN(n432) );
  NAND2_X1 U435 ( .A1(n431), .A2(n430), .ZN(n429) );
  INV_X1 U436 ( .A(n488), .ZN(n430) );
  INV_X1 U437 ( .A(G902), .ZN(n487) );
  XNOR2_X1 U438 ( .A(G113), .B(KEYINPUT87), .ZN(n438) );
  XNOR2_X1 U439 ( .A(n407), .B(G119), .ZN(n439) );
  XNOR2_X1 U440 ( .A(n416), .B(KEYINPUT93), .ZN(n415) );
  XNOR2_X1 U441 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n414) );
  INV_X1 U442 ( .A(n456), .ZN(n457) );
  XNOR2_X1 U443 ( .A(G122), .B(KEYINPUT9), .ZN(n518) );
  XOR2_X1 U444 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n519) );
  XNOR2_X1 U445 ( .A(G116), .B(G107), .ZN(n521) );
  INV_X1 U446 ( .A(G134), .ZN(n434) );
  XNOR2_X1 U447 ( .A(n423), .B(n422), .ZN(n525) );
  INV_X1 U448 ( .A(KEYINPUT8), .ZN(n422) );
  NAND2_X1 U449 ( .A1(n741), .A2(G234), .ZN(n423) );
  XOR2_X1 U450 ( .A(G137), .B(G140), .Z(n456) );
  INV_X1 U451 ( .A(KEYINPUT74), .ZN(n412) );
  INV_X1 U452 ( .A(KEYINPUT79), .ZN(n570) );
  XNOR2_X1 U453 ( .A(n515), .B(n380), .ZN(n517) );
  INV_X1 U454 ( .A(G475), .ZN(n380) );
  NAND2_X1 U455 ( .A1(n471), .A2(n470), .ZN(n573) );
  XNOR2_X1 U456 ( .A(n370), .B(n392), .ZN(n391) );
  INV_X1 U457 ( .A(KEYINPUT6), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n442), .B(n389), .ZN(n619) );
  XNOR2_X1 U459 ( .A(n390), .B(n437), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n415), .B(n414), .ZN(n437) );
  XNOR2_X1 U461 ( .A(n474), .B(n351), .ZN(n390) );
  NOR2_X1 U462 ( .A1(n420), .A2(n576), .ZN(n596) );
  NAND2_X1 U463 ( .A1(n405), .A2(n404), .ZN(n401) );
  INV_X1 U464 ( .A(KEYINPUT102), .ZN(n542) );
  INV_X1 U465 ( .A(KEYINPUT60), .ZN(n382) );
  INV_X1 U466 ( .A(G143), .ZN(n657) );
  AND2_X1 U467 ( .A1(n432), .A2(n427), .ZN(n348) );
  NOR2_X1 U468 ( .A1(n339), .A2(n545), .ZN(n349) );
  NOR2_X1 U469 ( .A1(n391), .A2(n419), .ZN(n350) );
  AND2_X1 U470 ( .A1(n508), .A2(G210), .ZN(n351) );
  AND2_X1 U471 ( .A1(n346), .A2(n391), .ZN(n352) );
  AND2_X1 U472 ( .A1(n555), .A2(n391), .ZN(n353) );
  AND2_X1 U473 ( .A1(n605), .A2(n628), .ZN(n354) );
  AND2_X1 U474 ( .A1(n428), .A2(n432), .ZN(n355) );
  XOR2_X1 U475 ( .A(n492), .B(KEYINPUT19), .Z(n356) );
  XNOR2_X1 U476 ( .A(n472), .B(KEYINPUT33), .ZN(n707) );
  NOR2_X1 U477 ( .A1(n561), .A2(n497), .ZN(n357) );
  XOR2_X1 U478 ( .A(n372), .B(n637), .Z(n359) );
  XOR2_X1 U479 ( .A(n619), .B(n618), .Z(n360) );
  XNOR2_X1 U480 ( .A(KEYINPUT122), .B(n613), .ZN(n361) );
  XOR2_X1 U481 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n363) );
  NAND2_X1 U482 ( .A1(n533), .A2(n552), .ZN(n697) );
  BUF_X1 U483 ( .A(n641), .Z(n717) );
  XNOR2_X1 U484 ( .A(n379), .B(n474), .ZN(n364) );
  BUF_X1 U485 ( .A(n640), .Z(n365) );
  XNOR2_X1 U486 ( .A(n379), .B(n474), .ZN(n728) );
  BUF_X1 U487 ( .A(n672), .Z(n366) );
  XNOR2_X1 U488 ( .A(n446), .B(n456), .ZN(n406) );
  XNOR2_X1 U489 ( .A(n442), .B(n406), .ZN(n644) );
  NOR2_X1 U490 ( .A1(n644), .A2(G902), .ZN(n374) );
  XNOR2_X1 U491 ( .A(n585), .B(KEYINPUT71), .ZN(n396) );
  NAND2_X1 U492 ( .A1(n396), .A2(n395), .ZN(n394) );
  BUF_X1 U493 ( .A(n587), .Z(n367) );
  BUF_X1 U494 ( .A(n660), .Z(n368) );
  XNOR2_X1 U495 ( .A(n387), .B(n570), .ZN(n660) );
  BUF_X1 U496 ( .A(n591), .Z(n369) );
  XNOR2_X2 U497 ( .A(n441), .B(n440), .ZN(n370) );
  BUF_X1 U498 ( .A(n344), .Z(n371) );
  XNOR2_X1 U499 ( .A(n728), .B(n484), .ZN(n638) );
  AND2_X1 U500 ( .A1(n679), .A2(n352), .ZN(n375) );
  XNOR2_X1 U501 ( .A(n408), .B(n362), .ZN(n378) );
  NAND2_X1 U502 ( .A1(n403), .A2(n530), .ZN(n376) );
  NAND2_X1 U503 ( .A1(n536), .A2(n679), .ZN(n541) );
  NAND2_X1 U504 ( .A1(n377), .A2(n631), .ZN(n544) );
  NOR2_X1 U505 ( .A1(n629), .A2(n640), .ZN(n377) );
  XNOR2_X1 U506 ( .A(n394), .B(KEYINPUT69), .ZN(n393) );
  NOR2_X2 U507 ( .A1(n747), .A2(n624), .ZN(n410) );
  XNOR2_X1 U508 ( .A(n507), .B(n506), .ZN(n514) );
  NOR2_X2 U509 ( .A1(n607), .A2(n606), .ZN(n612) );
  XNOR2_X1 U510 ( .A(n381), .B(n363), .ZN(G51) );
  NAND2_X1 U511 ( .A1(n386), .A2(n621), .ZN(n381) );
  XNOR2_X1 U512 ( .A(n383), .B(n382), .ZN(G60) );
  NAND2_X1 U513 ( .A1(n384), .A2(n621), .ZN(n383) );
  XNOR2_X1 U514 ( .A(n635), .B(n358), .ZN(n384) );
  XNOR2_X2 U515 ( .A(n385), .B(n443), .ZN(n475) );
  XNOR2_X1 U516 ( .A(n639), .B(n359), .ZN(n386) );
  NAND2_X1 U517 ( .A1(n393), .A2(n409), .ZN(n408) );
  NAND2_X1 U518 ( .A1(n421), .A2(n568), .ZN(n387) );
  XNOR2_X1 U519 ( .A(n388), .B(n477), .ZN(n478) );
  INV_X1 U520 ( .A(n669), .ZN(n395) );
  INV_X1 U521 ( .A(n502), .ZN(n398) );
  NAND2_X1 U522 ( .A1(n402), .A2(n401), .ZN(n532) );
  INV_X1 U523 ( .A(n707), .ZN(n405) );
  NAND2_X1 U524 ( .A1(n500), .A2(KEYINPUT34), .ZN(n403) );
  NAND2_X1 U525 ( .A1(n569), .A2(n357), .ZN(n499) );
  XNOR2_X1 U526 ( .A(n410), .B(KEYINPUT46), .ZN(n409) );
  XNOR2_X2 U527 ( .A(n411), .B(KEYINPUT39), .ZN(n599) );
  NAND2_X2 U528 ( .A1(n591), .A2(n694), .ZN(n411) );
  XNOR2_X2 U529 ( .A(n413), .B(n412), .ZN(n591) );
  NAND2_X1 U530 ( .A1(n579), .A2(n580), .ZN(n413) );
  NAND2_X1 U531 ( .A1(n418), .A2(n417), .ZN(n566) );
  INV_X1 U532 ( .A(n419), .ZN(n417) );
  INV_X1 U533 ( .A(n565), .ZN(n418) );
  INV_X1 U534 ( .A(n568), .ZN(n420) );
  NOR2_X2 U535 ( .A1(n660), .A2(n571), .ZN(n572) );
  NAND2_X1 U536 ( .A1(n343), .A2(n353), .ZN(n648) );
  XNOR2_X2 U537 ( .A(n535), .B(n424), .ZN(n536) );
  XNOR2_X1 U538 ( .A(n425), .B(n361), .ZN(n615) );
  NAND2_X1 U539 ( .A1(n617), .A2(G217), .ZN(n425) );
  INV_X1 U540 ( .A(KEYINPUT64), .ZN(n426) );
  INV_X1 U541 ( .A(n690), .ZN(n427) );
  XOR2_X1 U542 ( .A(n504), .B(n503), .Z(n433) );
  INV_X1 U543 ( .A(G110), .ZN(n449) );
  XNOR2_X1 U544 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n441), .B(n440), .ZN(n565) );
  BUF_X1 U547 ( .A(n610), .Z(n722) );
  XNOR2_X1 U548 ( .A(n475), .B(n445), .ZN(n446) );
  INV_X1 U549 ( .A(n721), .ZN(n621) );
  XOR2_X1 U550 ( .A(KEYINPUT73), .B(n436), .Z(n508) );
  XOR2_X1 U551 ( .A(G472), .B(KEYINPUT94), .Z(n440) );
  XNOR2_X2 U552 ( .A(G101), .B(KEYINPUT72), .ZN(n444) );
  NAND2_X1 U553 ( .A1(G227), .A2(n741), .ZN(n445) );
  XOR2_X1 U554 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n448) );
  XNOR2_X1 U555 ( .A(KEYINPUT70), .B(KEYINPUT77), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n448), .B(n447), .ZN(n452) );
  XNOR2_X1 U557 ( .A(G128), .B(G119), .ZN(n450) );
  XNOR2_X1 U558 ( .A(n452), .B(n451), .ZN(n454) );
  NAND2_X1 U559 ( .A1(n525), .A2(G221), .ZN(n453) );
  XNOR2_X1 U560 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X2 U561 ( .A(n455), .B(G146), .ZN(n481) );
  XNOR2_X1 U562 ( .A(n501), .B(n457), .ZN(n734) );
  XNOR2_X1 U563 ( .A(n458), .B(n734), .ZN(n613) );
  NAND2_X1 U564 ( .A1(n613), .A2(n487), .ZN(n466) );
  XOR2_X1 U565 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n462) );
  XNOR2_X2 U566 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n459) );
  XNOR2_X2 U567 ( .A(n459), .B(G902), .ZN(n606) );
  NAND2_X1 U568 ( .A1(n606), .A2(G234), .ZN(n460) );
  XNOR2_X2 U569 ( .A(KEYINPUT20), .B(n460), .ZN(n467) );
  NAND2_X1 U570 ( .A1(n467), .A2(G217), .ZN(n461) );
  XNOR2_X1 U571 ( .A(n462), .B(n461), .ZN(n464) );
  INV_X1 U572 ( .A(KEYINPUT90), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X2 U574 ( .A(n466), .B(n465), .ZN(n679) );
  INV_X1 U575 ( .A(n679), .ZN(n471) );
  NAND2_X1 U576 ( .A1(G221), .A2(n467), .ZN(n469) );
  XOR2_X1 U577 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n468) );
  XNOR2_X1 U578 ( .A(n469), .B(n468), .ZN(n678) );
  INV_X1 U579 ( .A(n678), .ZN(n470) );
  INV_X1 U580 ( .A(n573), .ZN(n681) );
  NAND2_X1 U581 ( .A1(n537), .A2(n681), .ZN(n545) );
  NAND2_X1 U582 ( .A1(n741), .A2(G224), .ZN(n476) );
  XNOR2_X1 U583 ( .A(n476), .B(KEYINPUT88), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U585 ( .A(n606), .ZN(n485) );
  NAND2_X1 U586 ( .A1(n487), .A2(n486), .ZN(n489) );
  NAND2_X1 U587 ( .A1(n489), .A2(G210), .ZN(n488) );
  NAND2_X1 U588 ( .A1(n489), .A2(G214), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n490), .B(KEYINPUT89), .ZN(n690) );
  INV_X1 U590 ( .A(KEYINPUT84), .ZN(n491) );
  INV_X1 U591 ( .A(KEYINPUT75), .ZN(n492) );
  NAND2_X1 U592 ( .A1(G234), .A2(G237), .ZN(n493) );
  XNOR2_X1 U593 ( .A(n493), .B(KEYINPUT14), .ZN(n677) );
  NOR2_X1 U594 ( .A1(G902), .A2(n741), .ZN(n495) );
  NOR2_X1 U595 ( .A1(G953), .A2(G952), .ZN(n494) );
  NOR2_X1 U596 ( .A1(n495), .A2(n494), .ZN(n496) );
  NAND2_X1 U597 ( .A1(n677), .A2(n496), .ZN(n561) );
  AND2_X1 U598 ( .A1(G953), .A2(G898), .ZN(n497) );
  INV_X1 U599 ( .A(KEYINPUT0), .ZN(n498) );
  XNOR2_X2 U600 ( .A(n499), .B(n498), .ZN(n550) );
  INV_X1 U601 ( .A(n550), .ZN(n500) );
  XOR2_X1 U602 ( .A(n501), .B(G140), .Z(n507) );
  XOR2_X1 U603 ( .A(n398), .B(G104), .Z(n505) );
  NAND2_X1 U604 ( .A1(G214), .A2(n508), .ZN(n510) );
  XOR2_X1 U605 ( .A(n510), .B(n509), .Z(n511) );
  XNOR2_X1 U606 ( .A(n512), .B(n511), .ZN(n513) );
  NOR2_X1 U607 ( .A1(G902), .A2(n634), .ZN(n515) );
  INV_X1 U608 ( .A(KEYINPUT13), .ZN(n516) );
  XNOR2_X1 U609 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U610 ( .A(n520), .B(KEYINPUT7), .Z(n522) );
  XNOR2_X1 U611 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U612 ( .A(n524), .B(n523), .Z(n527) );
  NAND2_X1 U613 ( .A1(G217), .A2(n525), .ZN(n526) );
  XNOR2_X1 U614 ( .A(n527), .B(n526), .ZN(n718) );
  NOR2_X1 U615 ( .A1(G902), .A2(n718), .ZN(n528) );
  XNOR2_X1 U616 ( .A(G478), .B(n528), .ZN(n552) );
  INV_X1 U617 ( .A(n552), .ZN(n529) );
  NAND2_X1 U618 ( .A1(n553), .A2(n529), .ZN(n582) );
  INV_X1 U619 ( .A(n582), .ZN(n530) );
  XNOR2_X1 U620 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n532), .B(n531), .ZN(n640) );
  INV_X1 U622 ( .A(n553), .ZN(n533) );
  NOR2_X1 U623 ( .A1(n697), .A2(n678), .ZN(n534) );
  NAND2_X1 U624 ( .A1(n550), .A2(n534), .ZN(n535) );
  INV_X1 U625 ( .A(n346), .ZN(n539) );
  NAND2_X1 U626 ( .A1(n339), .A2(n539), .ZN(n540) );
  XNOR2_X1 U627 ( .A(n543), .B(n542), .ZN(n631) );
  AND2_X1 U628 ( .A1(n550), .A2(n349), .ZN(n547) );
  XNOR2_X1 U629 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n546) );
  XNOR2_X1 U630 ( .A(n547), .B(n546), .ZN(n667) );
  INV_X1 U631 ( .A(n567), .ZN(n576) );
  OR2_X1 U632 ( .A1(n576), .A2(n573), .ZN(n548) );
  NOR2_X1 U633 ( .A1(n418), .A2(n548), .ZN(n549) );
  AND2_X1 U634 ( .A1(n550), .A2(n549), .ZN(n651) );
  NOR2_X1 U635 ( .A1(n667), .A2(n651), .ZN(n551) );
  XOR2_X1 U636 ( .A(KEYINPUT96), .B(n551), .Z(n554) );
  NOR2_X1 U637 ( .A1(n553), .A2(n552), .ZN(n666) );
  NOR2_X1 U638 ( .A1(n666), .A2(n663), .ZN(n571) );
  INV_X1 U639 ( .A(n571), .ZN(n691) );
  NAND2_X1 U640 ( .A1(n554), .A2(n691), .ZN(n556) );
  NOR2_X1 U641 ( .A1(n679), .A2(n346), .ZN(n555) );
  NAND2_X1 U642 ( .A1(n556), .A2(n648), .ZN(n557) );
  NOR2_X2 U643 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U644 ( .A(KEYINPUT45), .ZN(n559) );
  INV_X1 U645 ( .A(n561), .ZN(n563) );
  NAND2_X1 U646 ( .A1(G953), .A2(G900), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n563), .A2(n562), .ZN(n574) );
  NOR2_X1 U648 ( .A1(n678), .A2(n574), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n572), .B(KEYINPUT47), .ZN(n584) );
  OR2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n580) );
  XNOR2_X1 U652 ( .A(KEYINPUT30), .B(KEYINPUT104), .ZN(n578) );
  XNOR2_X1 U653 ( .A(n578), .B(n577), .ZN(n579) );
  NOR2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n369), .A2(n583), .ZN(n656) );
  NAND2_X1 U656 ( .A1(n584), .A2(n656), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n350), .B(KEYINPUT103), .ZN(n586) );
  INV_X1 U658 ( .A(n663), .ZN(n659) );
  NAND2_X1 U659 ( .A1(n602), .A2(n367), .ZN(n589) );
  XNOR2_X1 U660 ( .A(KEYINPUT83), .B(KEYINPUT36), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n581), .B(KEYINPUT38), .ZN(n694) );
  NAND2_X1 U663 ( .A1(n599), .A2(n663), .ZN(n593) );
  XNOR2_X1 U664 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n593), .B(n592), .ZN(n747) );
  NOR2_X1 U666 ( .A1(n697), .A2(n690), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n594), .A2(n694), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n708), .A2(n596), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n597) );
  XNOR2_X1 U670 ( .A(n598), .B(n597), .ZN(n624) );
  NAND2_X1 U671 ( .A1(n599), .A2(n666), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT107), .ZN(n745) );
  INV_X1 U673 ( .A(n745), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n690), .A2(n346), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(KEYINPUT43), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n604), .A2(n581), .ZN(n628) );
  NAND2_X1 U678 ( .A1(n344), .A2(KEYINPUT2), .ZN(n609) );
  INV_X1 U679 ( .A(KEYINPUT82), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n611), .A2(n722), .ZN(n676) );
  INV_X1 U682 ( .A(G952), .ZN(n614) );
  AND2_X1 U683 ( .A1(n614), .A2(G953), .ZN(n721) );
  NAND2_X1 U684 ( .A1(n615), .A2(n621), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n616), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U686 ( .A1(n617), .A2(G472), .ZN(n620) );
  XNOR2_X1 U687 ( .A(KEYINPUT85), .B(KEYINPUT62), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n620), .B(n360), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U690 ( .A(n623), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U691 ( .A(n624), .B(G137), .Z(G39) );
  INV_X1 U692 ( .A(n666), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n368), .A2(n625), .ZN(n627) );
  XNOR2_X1 U694 ( .A(G128), .B(KEYINPUT29), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n627), .B(n626), .ZN(G30) );
  XNOR2_X1 U696 ( .A(n628), .B(G140), .ZN(G42) );
  XOR2_X1 U697 ( .A(n629), .B(G119), .Z(G21) );
  XNOR2_X1 U698 ( .A(G110), .B(KEYINPUT110), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(G12) );
  XNOR2_X2 U700 ( .A(n345), .B(n426), .ZN(n641) );
  NAND2_X1 U701 ( .A1(n641), .A2(G475), .ZN(n635) );
  XNOR2_X1 U702 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n633) );
  NAND2_X1 U703 ( .A1(n641), .A2(G210), .ZN(n639) );
  XNOR2_X1 U704 ( .A(KEYINPUT80), .B(KEYINPUT54), .ZN(n636) );
  XOR2_X1 U705 ( .A(n636), .B(KEYINPUT55), .Z(n637) );
  XOR2_X1 U706 ( .A(G122), .B(n365), .Z(G24) );
  NAND2_X1 U707 ( .A1(n717), .A2(G469), .ZN(n646) );
  XNOR2_X1 U708 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT58), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U711 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n647), .A2(n721), .ZN(G54) );
  XNOR2_X1 U713 ( .A(G101), .B(n648), .ZN(G3) );
  NAND2_X1 U714 ( .A1(n651), .A2(n663), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n649), .B(KEYINPUT108), .ZN(n650) );
  XNOR2_X1 U716 ( .A(G104), .B(n650), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n653) );
  NAND2_X1 U718 ( .A1(n651), .A2(n666), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n653), .B(n652), .ZN(n655) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .Z(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(G9) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U723 ( .A(n658), .B(KEYINPUT111), .ZN(G45) );
  NOR2_X1 U724 ( .A1(n368), .A2(n659), .ZN(n661) );
  XOR2_X1 U725 ( .A(KEYINPUT112), .B(n661), .Z(n662) );
  XNOR2_X1 U726 ( .A(G146), .B(n662), .ZN(G48) );
  XOR2_X1 U727 ( .A(G113), .B(KEYINPUT113), .Z(n665) );
  NAND2_X1 U728 ( .A1(n667), .A2(n663), .ZN(n664) );
  XNOR2_X1 U729 ( .A(n665), .B(n664), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U731 ( .A(n668), .B(G116), .ZN(G18) );
  XNOR2_X1 U732 ( .A(n669), .B(KEYINPUT37), .ZN(n670) );
  XNOR2_X1 U733 ( .A(n670), .B(KEYINPUT114), .ZN(n671) );
  XNOR2_X1 U734 ( .A(G125), .B(n671), .ZN(G27) );
  XOR2_X1 U735 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n715) );
  INV_X1 U736 ( .A(n366), .ZN(n674) );
  XNOR2_X1 U737 ( .A(KEYINPUT81), .B(KEYINPUT2), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n712) );
  NAND2_X1 U740 ( .A1(G952), .A2(n677), .ZN(n705) );
  NAND2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n680), .B(KEYINPUT49), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n681), .A2(n346), .ZN(n682) );
  XOR2_X1 U744 ( .A(KEYINPUT50), .B(n682), .Z(n683) );
  NAND2_X1 U745 ( .A1(n339), .A2(n683), .ZN(n684) );
  NOR2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U747 ( .A1(n349), .A2(n686), .ZN(n687) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(n687), .Z(n689) );
  INV_X1 U749 ( .A(n708), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n702) );
  NAND2_X1 U751 ( .A1(n691), .A2(n427), .ZN(n693) );
  INV_X1 U752 ( .A(n694), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n699) );
  NOR2_X1 U754 ( .A1(n694), .A2(n427), .ZN(n695) );
  XNOR2_X1 U755 ( .A(n695), .B(KEYINPUT116), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n700), .A2(n707), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U760 ( .A(n703), .B(KEYINPUT52), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U762 ( .A(KEYINPUT117), .B(n706), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n405), .A2(n708), .ZN(n709) );
  NAND2_X1 U764 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n713), .A2(n741), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U768 ( .A(KEYINPUT118), .B(n716), .Z(G75) );
  NAND2_X1 U769 ( .A1(n717), .A2(G478), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n720), .A2(n721), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n722), .A2(n741), .ZN(n727) );
  NAND2_X1 U773 ( .A1(G224), .A2(G953), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n724), .ZN(n725) );
  NAND2_X1 U776 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U777 ( .A1(n727), .A2(n726), .ZN(n732) );
  INV_X1 U778 ( .A(n364), .ZN(n730) );
  NOR2_X1 U779 ( .A1(G898), .A2(n741), .ZN(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT125), .B(n733), .Z(G69) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(n739) );
  XOR2_X1 U784 ( .A(G227), .B(n739), .Z(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U786 ( .A1(G953), .A2(n737), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(KEYINPUT126), .ZN(n744) );
  XNOR2_X1 U788 ( .A(n371), .B(n739), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U790 ( .A1(n744), .A2(n743), .ZN(G72) );
  XNOR2_X1 U791 ( .A(G134), .B(n745), .ZN(n746) );
  XNOR2_X1 U792 ( .A(n746), .B(KEYINPUT115), .ZN(G36) );
  BUF_X1 U793 ( .A(n747), .Z(n748) );
  XOR2_X1 U794 ( .A(G131), .B(n748), .Z(G33) );
endmodule

