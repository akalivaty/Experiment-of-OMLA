//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n204));
  INV_X1    g0004(.A(G58), .ZN(new_n205));
  INV_X1    g0005(.A(G232), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n203), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n203), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n205), .A2(new_n207), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n217), .A2(new_n218), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n217), .B2(new_n218), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n214), .A2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n206), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G68), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(KEYINPUT13), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  AND2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  OAI211_X1 g0047(.A(G226), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT72), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(KEYINPUT72), .A3(G226), .A4(new_n245), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G97), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n250), .A2(new_n252), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT73), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(KEYINPUT73), .A3(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT66), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n219), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n262), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n266), .A2(new_n262), .A3(new_n269), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT67), .B(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n268), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n256), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n271), .A2(new_n272), .B1(G238), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n244), .B1(new_n261), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n255), .A2(KEYINPUT73), .A3(new_n256), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT73), .B1(new_n255), .B2(new_n256), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n244), .B(new_n276), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(G169), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n277), .A2(new_n281), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n282), .A2(KEYINPUT14), .B1(new_n283), .B2(G179), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n282), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT13), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(new_n280), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT14), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n284), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n219), .B1(new_n203), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G50), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n297), .A2(new_n298), .B1(new_n220), .B2(G68), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n220), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G77), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  INV_X1    g0104(.A(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT67), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G1), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n306), .A2(new_n308), .A3(G13), .A4(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n273), .A2(new_n311), .A3(G13), .A4(G20), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT12), .A3(new_n207), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n304), .B(new_n314), .C1(KEYINPUT12), .C2(new_n313), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n273), .A2(G20), .ZN(new_n317));
  INV_X1    g0117(.A(new_n295), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n207), .B1(new_n319), .B2(KEYINPUT12), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n293), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n289), .A2(new_n280), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(G200), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n283), .A2(G190), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n317), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n316), .A2(new_n318), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n316), .A2(new_n330), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT78), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  INV_X1    g0139(.A(new_n337), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT69), .B1(new_n316), .B2(new_n318), .ZN(new_n341));
  AOI211_X1 g0141(.A(new_n333), .B(new_n295), .C1(new_n310), .C2(new_n312), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n339), .B(new_n340), .C1(new_n343), .C2(new_n331), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  AND3_X1   g0145(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT75), .B1(G58), .B2(G68), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n220), .B1(new_n348), .B2(new_n222), .ZN(new_n349));
  INV_X1    g0149(.A(G159), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n297), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n246), .A2(new_n247), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n353), .B2(new_n220), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NOR4_X1   g0155(.A1(new_n246), .A2(new_n247), .A3(new_n355), .A4(G20), .ZN(new_n356));
  OAI21_X1  g0156(.A(G68), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n222), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(new_n351), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT76), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n352), .A2(new_n357), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n357), .A4(new_n365), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n295), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n338), .A2(new_n344), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n251), .A2(G226), .ZN(new_n372));
  INV_X1    g0172(.A(G87), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n372), .A2(new_n245), .B1(new_n294), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n245), .A2(G223), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n353), .B2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n251), .A2(KEYINPUT79), .A3(G223), .A4(new_n245), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n256), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT80), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT80), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n377), .A2(new_n378), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n382), .B(new_n256), .C1(new_n383), .C2(new_n374), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n275), .A2(G232), .ZN(new_n385));
  INV_X1    g0185(.A(G179), .ZN(new_n386));
  INV_X1    g0186(.A(new_n272), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n270), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n381), .A2(new_n384), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n379), .A2(new_n380), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n271), .A2(new_n272), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n385), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n287), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n371), .A2(new_n395), .A3(KEYINPUT18), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT18), .B1(new_n371), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT81), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n371), .A2(new_n395), .A3(KEYINPUT81), .A4(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n338), .A2(new_n344), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G200), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n391), .B2(new_n393), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n381), .A2(new_n384), .ZN(new_n406));
  INV_X1    g0206(.A(G190), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n392), .A2(new_n407), .A3(new_n385), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n370), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT17), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n403), .A2(new_n412), .A3(new_n370), .A4(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n401), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT70), .B1(new_n353), .B2(new_n206), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT70), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n251), .A2(new_n418), .A3(G232), .A4(new_n245), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n417), .B(new_n419), .C1(new_n420), .C2(new_n251), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n251), .A2(G238), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n245), .B1(new_n422), .B2(new_n418), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n256), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n271), .A2(new_n272), .B1(G244), .B2(new_n275), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n386), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n319), .A2(new_n301), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n300), .B1(new_n220), .B2(new_n301), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n329), .A2(new_n297), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n295), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G77), .B2(new_n316), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n426), .A2(new_n287), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n428), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n427), .A2(new_n404), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n426), .B2(new_n407), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n245), .A2(G222), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G223), .A2(G1698), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n251), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n256), .C1(G77), .C2(new_n251), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n275), .A2(G226), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n392), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G169), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n386), .B2(new_n447), .ZN(new_n449));
  OAI211_X1 g0249(.A(G50), .B(new_n317), .C1(new_n341), .C2(new_n342), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n296), .A2(G150), .ZN(new_n451));
  NOR3_X1   g0251(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n452));
  OAI221_X1 g0252(.A(new_n451), .B1(new_n452), .B2(new_n220), .C1(new_n329), .C2(new_n300), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n313), .A2(new_n298), .B1(new_n295), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n455), .A2(KEYINPUT9), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n455), .A2(KEYINPUT9), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT71), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n447), .A2(new_n404), .ZN(new_n461));
  AOI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(G190), .C2(new_n447), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT10), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT10), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n459), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n441), .B(new_n456), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n328), .A2(new_n416), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT82), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n220), .B1(new_n471), .B2(G33), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G20), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n295), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n469), .A2(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n469), .A2(KEYINPUT82), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n295), .A2(new_n476), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n313), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n273), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n316), .A2(G116), .A3(new_n318), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(KEYINPUT86), .A2(G303), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT86), .A2(G303), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n353), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n245), .A2(G257), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G264), .A2(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n251), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n494), .A3(new_n256), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT87), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT87), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(new_n494), .A3(new_n497), .A4(new_n256), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT5), .B(G41), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n306), .A2(new_n308), .A3(G45), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n380), .B(G270), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n502), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n266), .A3(new_n500), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND4_X1   g0306(.A1(G179), .A2(new_n488), .A3(new_n499), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n287), .B1(new_n499), .B2(new_n506), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n488), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT21), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n511), .A3(new_n488), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n507), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n499), .A2(new_n506), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G200), .ZN(new_n515));
  INV_X1    g0315(.A(new_n488), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n407), .C2(new_n514), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n245), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n470), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n256), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n380), .B(G257), .C1(new_n501), .C2(new_n502), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(new_n505), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n287), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n531), .A2(new_n471), .A3(G107), .ZN(new_n532));
  XNOR2_X1  g0332(.A(G97), .B(G107), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n534), .A2(new_n220), .B1(new_n301), .B2(new_n297), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n355), .B1(new_n251), .B2(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n353), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n420), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n295), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n316), .A2(G97), .A3(new_n318), .A4(new_n486), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n313), .A2(new_n471), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n527), .A2(new_n505), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT83), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n527), .A2(new_n505), .A3(KEYINPUT83), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n526), .A3(new_n386), .A4(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n530), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n543), .A2(new_n544), .B1(new_n525), .B2(new_n256), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G200), .ZN(new_n551));
  INV_X1    g0351(.A(new_n542), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT84), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n526), .A2(new_n528), .A3(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n540), .A3(new_n541), .A4(new_n539), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n404), .B1(new_n549), .B2(new_n546), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT84), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n548), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  AND4_X1   g0359(.A1(G107), .A2(new_n316), .A3(new_n318), .A4(new_n486), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n220), .B(G87), .C1(new_n246), .C2(new_n247), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n251), .A2(new_n563), .A3(new_n220), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT88), .B1(new_n566), .B2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT88), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(new_n220), .A3(G33), .A4(G116), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT23), .B1(new_n220), .B2(G107), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n420), .A3(G20), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n567), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n318), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n562), .B2(new_n564), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT24), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n560), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT25), .A4(new_n420), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT25), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n316), .B2(G107), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G250), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G257), .A2(G1698), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n589), .C1(new_n353), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n256), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n380), .B(G264), .C1(new_n501), .C2(new_n502), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n505), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G169), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G179), .ZN(new_n597));
  INV_X1    g0397(.A(new_n505), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n587), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n504), .A2(new_n263), .ZN(new_n602));
  INV_X1    g0402(.A(G250), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n502), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n380), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n566), .B1(new_n422), .B2(G1698), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(G1698), .C1(new_n246), .C2(new_n247), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n386), .B(new_n605), .C1(new_n610), .C2(new_n380), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n310), .A2(new_n312), .A3(new_n430), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n251), .A2(new_n220), .A3(G68), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n373), .A2(new_n471), .A3(new_n420), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n253), .A2(new_n220), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT19), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n300), .B2(new_n471), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n295), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n316), .A2(new_n318), .A3(new_n486), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n612), .B(new_n620), .C1(new_n621), .C2(new_n430), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n607), .B(KEYINPUT85), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n353), .A2(new_n208), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n245), .B1(G33), .B2(G116), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n380), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n605), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n611), .B(new_n622), .C1(new_n628), .C2(G169), .ZN(new_n629));
  OAI21_X1  g0429(.A(G200), .B1(new_n626), .B2(new_n627), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n316), .A2(G87), .A3(new_n318), .A4(new_n486), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n620), .A2(new_n612), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(G190), .B(new_n605), .C1(new_n610), .C2(new_n380), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n594), .A2(G200), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n596), .A2(G190), .A3(new_n505), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n580), .A2(new_n586), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n601), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n468), .A2(new_n519), .A3(new_n559), .A4(new_n642), .ZN(G372));
  AND3_X1   g0443(.A1(new_n371), .A2(new_n395), .A3(KEYINPUT18), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT92), .B1(new_n644), .B2(new_n397), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n371), .A2(new_n395), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n396), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n438), .B1(new_n325), .B2(new_n326), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n293), .B2(new_n322), .ZN(new_n653));
  INV_X1    g0453(.A(new_n414), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n464), .A2(new_n466), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n456), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(KEYINPUT93), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n629), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT90), .B1(new_n632), .B2(new_n633), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT90), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n631), .A2(new_n666), .A3(new_n612), .A4(new_n620), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n630), .A3(new_n635), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n640), .A2(new_n668), .A3(new_n629), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n513), .B2(new_n600), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n664), .B1(new_n670), .B2(new_n559), .ZN(new_n671));
  INV_X1    g0471(.A(new_n637), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n548), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n548), .A2(new_n668), .A3(new_n629), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n548), .A2(new_n636), .A3(new_n629), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n676), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n673), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n671), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n468), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n663), .A2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(new_n513), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n220), .A2(G13), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n273), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  OAI21_X1  g0487(.A(G213), .B1(new_n686), .B2(KEYINPUT27), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n516), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n518), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n601), .A2(new_n641), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n587), .A2(new_n691), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n600), .B2(new_n692), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n513), .A2(new_n691), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n698), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n601), .A2(new_n692), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n702), .A2(new_n707), .ZN(G399));
  OR2_X1    g0508(.A1(new_n614), .A2(G116), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  INV_X1    g0510(.A(new_n215), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G1), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n710), .A2(new_n714), .B1(new_n223), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(G330), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n596), .A2(G179), .ZN(new_n718));
  INV_X1    g0518(.A(new_n514), .ZN(new_n719));
  INV_X1    g0519(.A(new_n529), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(new_n628), .ZN(new_n721));
  XNOR2_X1  g0521(.A(KEYINPUT95), .B(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n628), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n594), .A2(new_n386), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n514), .A3(new_n550), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT96), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n721), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n723), .A2(KEYINPUT96), .A3(new_n726), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n692), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n723), .A3(new_n726), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n691), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n733), .A2(new_n735), .B1(new_n737), .B2(new_n734), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n519), .A2(new_n559), .A3(new_n642), .A4(new_n692), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n717), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n681), .A2(new_n692), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n555), .A2(new_n558), .ZN(new_n744));
  INV_X1    g0544(.A(new_n548), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT97), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n559), .A2(KEYINPUT97), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(new_n670), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n629), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(KEYINPUT26), .B2(new_n675), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n691), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT29), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n740), .B1(new_n743), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n716), .B1(new_n755), .B2(G1), .ZN(G364));
  AOI21_X1  g0556(.A(new_n305), .B1(new_n685), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n712), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n697), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n695), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n219), .B1(G20), .B2(new_n287), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n220), .A2(new_n407), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n386), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n220), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n766), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n767), .A2(new_n205), .B1(new_n769), .B2(new_n301), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n404), .A2(G179), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n353), .B(new_n770), .C1(G87), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n220), .B1(new_n775), .B2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n471), .ZN(new_n777));
  NAND3_X1  g0577(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n407), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n298), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(G190), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n777), .B(new_n781), .C1(G68), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n768), .A2(new_n775), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n350), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n771), .A2(new_n768), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT98), .Z(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G107), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n774), .A2(new_n783), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n353), .B1(new_n772), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G326), .B2(new_n779), .ZN(new_n794));
  INV_X1    g0594(.A(new_n776), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n795), .A2(G294), .B1(new_n782), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n767), .A2(new_n798), .B1(new_n769), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n784), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G329), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n791), .A2(new_n794), .A3(new_n797), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n764), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n239), .A2(G45), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n711), .A2(new_n251), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(G45), .C2(new_n223), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n711), .A2(new_n353), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G355), .B1(new_n475), .B2(new_n711), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n763), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n762), .B(new_n804), .C1(new_n810), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n813), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n695), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n761), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n438), .A2(new_n691), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n440), .A2(new_n439), .B1(new_n435), .B2(new_n692), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n438), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n741), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n824), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n681), .A2(new_n692), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n740), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n713), .B2(new_n757), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n740), .A2(new_n825), .A3(new_n827), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n763), .A2(new_n811), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n762), .B1(new_n301), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n353), .B1(new_n772), .B2(new_n420), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT99), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n780), .A2(new_n792), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n777), .B(new_n836), .C1(G283), .C2(new_n782), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n788), .A2(G87), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n767), .A2(new_n839), .B1(new_n784), .B2(new_n799), .ZN(new_n840));
  INV_X1    g0640(.A(new_n769), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(G116), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g0642(.A1(new_n835), .A2(new_n837), .A3(new_n838), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n251), .B1(new_n784), .B2(new_n844), .C1(new_n298), .C2(new_n772), .ZN(new_n845));
  INV_X1    g0645(.A(new_n788), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n207), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(G58), .C2(new_n795), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT100), .ZN(new_n849));
  INV_X1    g0649(.A(new_n767), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n850), .B1(new_n841), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  INV_X1    g0652(.A(G150), .ZN(new_n853));
  INV_X1    g0653(.A(new_n782), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n851), .B1(new_n780), .B2(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n843), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n833), .B1(new_n857), .B2(new_n764), .C1(new_n812), .C2(new_n826), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n831), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  INV_X1    g0660(.A(new_n534), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n861), .A2(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(KEYINPUT35), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(G116), .A3(new_n221), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  NAND3_X1  g0665(.A1(new_n224), .A2(G77), .A3(new_n348), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT101), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n866), .A2(KEYINPUT101), .B1(new_n298), .B2(G68), .ZN(new_n868));
  AOI211_X1 g0668(.A(G13), .B(new_n273), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n369), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT104), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n357), .A2(new_n365), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT76), .B1(new_n363), .B2(new_n364), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n352), .A2(KEYINPUT104), .A3(new_n357), .A4(new_n365), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n367), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n295), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n871), .B1(new_n878), .B2(KEYINPUT105), .ZN(new_n879));
  INV_X1    g0679(.A(new_n367), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n366), .B2(new_n872), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n318), .B1(new_n881), .B2(new_n876), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n402), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n689), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n415), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n395), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n410), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  XOR2_X1   g0690(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n891));
  INV_X1    g0691(.A(new_n689), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n371), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n410), .A2(new_n646), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n887), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(new_n894), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n369), .B1(new_n882), .B2(new_n883), .ZN(new_n899));
  AOI211_X1 g0699(.A(KEYINPUT105), .B(new_n318), .C1(new_n881), .C2(new_n876), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n403), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n892), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n395), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n410), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n898), .B1(new_n904), .B2(KEYINPUT37), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n401), .B2(new_n414), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n321), .A2(new_n692), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n290), .A2(new_n291), .B1(new_n324), .B2(new_n386), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT74), .B1(new_n282), .B2(KEYINPUT14), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n290), .A2(new_n286), .A3(new_n291), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n327), .B(new_n910), .C1(new_n914), .C2(new_n321), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT103), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n293), .A2(new_n909), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n737), .A2(new_n734), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n739), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n923), .A2(new_n826), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n908), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n915), .A2(new_n917), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT103), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n893), .B1(new_n651), .B2(new_n414), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n410), .A2(new_n646), .A3(new_n893), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(new_n891), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n897), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n926), .B1(new_n935), .B2(new_n896), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n925), .A2(new_n926), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n468), .A2(new_n923), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT107), .ZN(new_n940));
  OAI21_X1  g0740(.A(G330), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n938), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n323), .A2(new_n691), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n935), .A2(new_n896), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT102), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n691), .B(new_n824), .C1(new_n671), .C2(new_n680), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n820), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n827), .A2(KEYINPUT102), .A3(new_n821), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n908), .A3(new_n920), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n645), .A2(new_n650), .A3(new_n689), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n468), .A2(new_n743), .A3(new_n754), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n663), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n942), .A2(new_n960), .B1(new_n273), .B2(new_n685), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n942), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n870), .B1(new_n961), .B2(new_n962), .ZN(G367));
  OAI211_X1 g0763(.A(new_n748), .B(new_n749), .C1(new_n552), .C2(new_n692), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n548), .A2(new_n691), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT109), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n964), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n704), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  INV_X1    g0773(.A(new_n970), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n745), .B1(new_n974), .B2(new_n600), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n692), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n665), .A2(new_n667), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n691), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n629), .A3(new_n668), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n629), .B2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT108), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n982), .B2(new_n981), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n985), .B1(new_n976), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n702), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n970), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n990), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n985), .B(new_n992), .C1(new_n976), .C2(new_n987), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n712), .B(KEYINPUT41), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n970), .A2(new_n707), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT45), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n967), .A2(new_n706), .A3(new_n969), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n1002), .A3(new_n702), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n704), .B1(new_n701), .B2(new_n703), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n697), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n989), .B1(new_n996), .B2(new_n1001), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n755), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n994), .B1(new_n1007), .B2(new_n755), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n991), .B(new_n993), .C1(new_n1008), .C2(new_n758), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n814), .B1(new_n215), .B2(new_n430), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n234), .B2(new_n806), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n772), .A2(new_n475), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(KEYINPUT46), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G107), .B2(new_n795), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1012), .A2(KEYINPUT46), .B1(G311), .B2(new_n779), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n489), .A2(new_n490), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(G283), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1017), .A2(new_n767), .B1(new_n769), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G317), .B2(new_n801), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n353), .B1(new_n787), .B2(new_n471), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G294), .B2(new_n782), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1014), .A2(new_n1015), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n776), .A2(new_n207), .ZN(new_n1024));
  INV_X1    g0824(.A(G143), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n780), .A2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(G159), .C2(new_n782), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n841), .B1(new_n801), .B2(G137), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G58), .A2(new_n773), .B1(new_n850), .B2(G150), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n251), .B1(new_n787), .B2(new_n301), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT110), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1023), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n762), .B(new_n1011), .C1(new_n1034), .C2(new_n763), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n981), .B2(new_n816), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1009), .A2(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n1005), .A2(new_n758), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n701), .A2(new_n816), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n788), .A2(G97), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n776), .A2(new_n430), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n353), .B(new_n1041), .C1(G50), .C2(new_n850), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n330), .A2(new_n782), .B1(G159), .B2(new_n779), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n769), .A2(new_n207), .B1(new_n784), .B2(new_n853), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G77), .B2(new_n773), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n251), .B1(new_n801), .B2(G326), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n772), .A2(new_n839), .B1(new_n776), .B2(new_n1018), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G317), .A2(new_n850), .B1(new_n841), .B2(new_n1016), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n780), .B2(new_n798), .C1(new_n799), .C2(new_n854), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1047), .B1(new_n475), .B2(new_n787), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1046), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n764), .B1(new_n1057), .B2(KEYINPUT113), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(KEYINPUT113), .B2(new_n1057), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n710), .A2(new_n808), .B1(new_n420), .B2(new_n711), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n710), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT111), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT111), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n329), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  AOI21_X1  g0865(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(new_n806), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT112), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n231), .A2(G45), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1068), .B2(KEYINPUT112), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1060), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n762), .B1(new_n1072), .B2(new_n814), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1059), .A2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n755), .A2(new_n1005), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n755), .A2(new_n1005), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n712), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1038), .B1(new_n1039), .B2(new_n1074), .C1(new_n1078), .C2(new_n1079), .ZN(G393));
  NAND3_X1  g0880(.A1(new_n1003), .A2(new_n758), .A3(new_n1006), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n806), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n814), .B1(new_n471), .B2(new_n215), .C1(new_n242), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n759), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n769), .A2(new_n329), .B1(new_n784), .B2(new_n1025), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n353), .B(new_n1085), .C1(G68), .C2(new_n773), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n776), .A2(new_n301), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n782), .B2(G50), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n838), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n850), .A2(G159), .B1(G150), .B2(new_n779), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n251), .B1(new_n773), .B2(G283), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G294), .A2(new_n841), .B1(new_n801), .B2(G322), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n795), .A2(G116), .B1(new_n1016), .B2(new_n782), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n789), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n850), .A2(G311), .B1(G317), .B2(new_n779), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1089), .A2(new_n1091), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1084), .B1(new_n1098), .B2(new_n763), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n970), .B2(new_n816), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1081), .A2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1007), .A2(new_n712), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1077), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  NAND3_X1  g0906(.A1(new_n923), .A2(G330), .A3(new_n826), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n918), .B2(new_n919), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n717), .B(new_n824), .C1(new_n738), .C2(new_n739), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n920), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n823), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n691), .B(new_n1113), .C1(new_n750), .C2(new_n752), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT115), .B1(new_n1114), .B2(new_n820), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n753), .A2(new_n823), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT115), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n821), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(KEYINPUT116), .B(new_n1107), .C1(new_n918), .C2(new_n919), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1110), .A2(new_n1112), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n920), .A2(new_n1111), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n918), .A2(new_n1107), .A3(new_n919), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n953), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n468), .A2(G330), .A3(new_n923), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT93), .B1(new_n657), .B2(new_n658), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n660), .B(new_n456), .C1(new_n655), .C2(new_n656), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n958), .B(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1123), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n946), .B1(new_n896), .B2(new_n907), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n935), .A2(new_n896), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n946), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n950), .A2(new_n949), .A3(new_n820), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT102), .B1(new_n827), .B2(new_n821), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n928), .A2(new_n929), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n944), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n943), .B1(new_n935), .B2(new_n896), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1119), .B2(new_n1139), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1132), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n945), .A2(new_n947), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n943), .B1(new_n953), .B2(new_n920), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1143), .B(new_n1112), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1131), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1123), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1129), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1147), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n712), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n758), .A3(new_n1147), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n769), .A2(new_n1156), .B1(new_n776), .B2(new_n350), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G137), .B2(new_n782), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT117), .Z(new_n1159));
  NOR2_X1   g0959(.A1(new_n772), .A2(new_n853), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n353), .B1(new_n801), .B2(G125), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n298), .B2(new_n787), .C1(new_n844), .C2(new_n767), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G128), .B2(new_n779), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n847), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n251), .B(new_n1087), .C1(G87), .C2(new_n773), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G107), .A2(new_n782), .B1(new_n779), .B2(G283), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n767), .A2(new_n475), .B1(new_n769), .B2(new_n471), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G294), .B2(new_n801), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n764), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n762), .B(new_n1172), .C1(new_n329), .C2(new_n832), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1145), .B2(new_n812), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1155), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1154), .A2(new_n1175), .ZN(G378));
  AND2_X1   g0976(.A1(new_n896), .A2(new_n907), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n926), .B1(new_n1177), .B2(new_n930), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n931), .A2(new_n936), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(G330), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n656), .B2(new_n658), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n456), .B(new_n1181), .C1(new_n464), .C2(new_n466), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n689), .B1(new_n450), .B2(new_n454), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OR3_X1    g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1180), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n937), .A2(G330), .A3(new_n1189), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n957), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n948), .A2(new_n956), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1189), .B1(new_n937), .B2(G330), .ZN(new_n1195));
  AND4_X1   g0995(.A1(G330), .A2(new_n1178), .A3(new_n1179), .A4(new_n1189), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1193), .A2(new_n1197), .B1(new_n1153), .B2(new_n1130), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n712), .B1(new_n1198), .B2(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1193), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1153), .A2(new_n1130), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1200), .A2(KEYINPUT57), .A3(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n832), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n759), .B1(G50), .B2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n767), .A2(new_n420), .B1(new_n784), .B2(new_n1018), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n430), .A2(new_n769), .B1(new_n787), .B2(new_n205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n267), .B(new_n353), .C1(new_n772), .C2(new_n301), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1207), .C1(KEYINPUT118), .C2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n780), .A2(new_n475), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1024), .B(new_n1210), .C1(G97), .C2(new_n782), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(KEYINPUT118), .C2(new_n1208), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT58), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n246), .A2(G41), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1212), .A2(new_n1213), .B1(new_n298), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1156), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n773), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT119), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n767), .A2(new_n1219), .B1(new_n769), .B2(new_n852), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G132), .B2(new_n782), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n795), .A2(G150), .B1(G125), .B2(new_n779), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1218), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n294), .B(new_n267), .C1(new_n787), .C2(new_n350), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G124), .B2(new_n801), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1215), .B1(new_n1213), .B2(new_n1212), .C1(new_n1224), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1205), .B1(new_n1229), .B2(new_n763), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1189), .B2(new_n812), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT120), .Z(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1200), .B2(new_n758), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1203), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G375));
  INV_X1    g1035(.A(new_n994), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1121), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1131), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n251), .B1(new_n788), .B2(G77), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT121), .Z(new_n1240));
  AOI21_X1  g1040(.A(new_n1041), .B1(new_n779), .B2(G294), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G283), .A2(new_n850), .B1(new_n841), .B2(G107), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G97), .A2(new_n773), .B1(new_n801), .B2(G303), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n782), .A2(G116), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n772), .A2(new_n350), .B1(new_n784), .B2(new_n1219), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT122), .Z(new_n1248));
  AOI22_X1  g1048(.A1(new_n1216), .A2(new_n782), .B1(G132), .B2(new_n779), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n298), .B2(new_n776), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n251), .B1(new_n787), .B2(new_n205), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n767), .A2(new_n852), .B1(new_n769), .B2(new_n853), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1248), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n763), .B1(new_n1246), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1254), .B(new_n759), .C1(G68), .C2(new_n1204), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1139), .B2(new_n811), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1125), .B2(new_n758), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(new_n1257), .ZN(G381));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G378), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1154), .A2(new_n1175), .A3(KEYINPUT123), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1009), .A2(new_n1105), .A3(new_n1036), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1234), .A2(new_n1263), .A3(new_n1265), .A4(new_n1266), .ZN(G407));
  NAND2_X1  g1067(.A1(new_n690), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1234), .A2(new_n1263), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  AOI21_X1  g1071(.A(new_n1105), .B1(new_n1009), .B2(new_n1036), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(G393), .B(new_n818), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1264), .A3(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1265), .B2(new_n1272), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT124), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1191), .A2(new_n1192), .A3(new_n957), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n957), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1197), .A2(KEYINPUT124), .A3(new_n1193), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1283), .A2(new_n758), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1200), .A2(new_n1236), .A3(new_n1201), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1232), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1260), .B(new_n1261), .C1(new_n1285), .C2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1233), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1237), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1237), .A2(new_n1292), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n712), .A3(new_n1131), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1257), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n859), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(G384), .A3(new_n1257), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1291), .A2(new_n1268), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1278), .B1(new_n1279), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1291), .A2(new_n1268), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1269), .A2(G2897), .ZN(new_n1304));
  XOR2_X1   g1104(.A(new_n1304), .B(KEYINPUT125), .Z(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1299), .B(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1303), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1301), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(KEYINPUT63), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1279), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1302), .B(new_n1308), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1269), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1314), .A2(KEYINPUT62), .A3(new_n1300), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT62), .B1(new_n1314), .B2(new_n1300), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1308), .B(KEYINPUT127), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1278), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1301), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1314), .A2(KEYINPUT62), .A3(new_n1300), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT127), .B1(new_n1322), .B2(new_n1308), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1313), .B1(new_n1318), .B2(new_n1323), .ZN(G405));
  OAI21_X1  g1124(.A(new_n1290), .B1(new_n1234), .B2(new_n1262), .ZN(new_n1325));
  OR2_X1    g1125(.A1(new_n1325), .A2(new_n1300), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1300), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1278), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1277), .A3(new_n1276), .A4(new_n1327), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(G402));
endmodule


