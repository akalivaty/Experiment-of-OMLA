//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n223), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n222), .A2(new_n225), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n229), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT64), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G222), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n253), .B(new_n255), .C1(new_n256), .C2(new_n254), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n250), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n257), .B(new_n260), .C1(G77), .C2(new_n253), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n259), .A2(new_n262), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n261), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G190), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(new_n273), .B1(G200), .B2(new_n268), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n203), .A2(G20), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT65), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(new_n250), .B2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n219), .A2(KEYINPUT65), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n275), .B1(new_n276), .B2(new_n278), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n224), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n284), .A2(new_n286), .B1(new_n202), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n285), .A2(new_n224), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n218), .A2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n202), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g0093(.A(new_n293), .B(KEYINPUT9), .Z(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n274), .A2(KEYINPUT10), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(new_n273), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n271), .B1(new_n299), .B2(new_n269), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n268), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT66), .B(G179), .Z(new_n304));
  OAI211_X1 g0104(.A(new_n293), .B(new_n303), .C1(new_n304), .C2(new_n268), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n296), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT16), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n251), .A2(new_n219), .A3(new_n252), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n252), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n214), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G58), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n214), .ZN(new_n314));
  OAI21_X1  g0114(.A(G20), .B1(new_n314), .B2(new_n201), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n277), .A2(G159), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n307), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n321), .B2(new_n219), .ZN(new_n322));
  INV_X1    g0122(.A(new_n311), .ZN(new_n323));
  OAI21_X1  g0123(.A(G68), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n317), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n326), .A3(new_n286), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n256), .A2(new_n254), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n213), .A2(G1698), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(new_n319), .C2(new_n320), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G87), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n260), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n259), .A2(G232), .A3(new_n262), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .A4(new_n265), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n259), .B1(new_n330), .B2(new_n331), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n338), .A2(new_n334), .A3(new_n264), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n339), .B2(G200), .ZN(new_n340));
  INV_X1    g0140(.A(new_n283), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n292), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n283), .A2(new_n287), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n342), .A2(KEYINPUT75), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT75), .B1(new_n342), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n327), .A2(new_n340), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT78), .A3(KEYINPUT17), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n327), .A2(new_n340), .A3(KEYINPUT78), .A4(new_n346), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n327), .A2(new_n346), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n333), .A2(new_n335), .A3(new_n265), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G169), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n339), .A2(new_n304), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT77), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n327), .A2(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT18), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT76), .ZN(new_n365));
  AND4_X1   g0165(.A1(new_n365), .A2(new_n353), .A3(KEYINPUT18), .A4(new_n357), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n361), .B2(KEYINPUT18), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n352), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n306), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  OAI211_X1 g0171(.A(G232), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT71), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n253), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  OAI211_X1 g0177(.A(G226), .B(new_n254), .C1(new_n319), .C2(new_n320), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n264), .B1(new_n379), .B2(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n259), .A2(new_n262), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n215), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n371), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n378), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n374), .B2(new_n375), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n259), .B1(new_n386), .B2(new_n377), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n387), .A2(KEYINPUT13), .A3(new_n382), .A4(new_n264), .ZN(new_n388));
  OAI21_X1  g0188(.A(G169), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT14), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT72), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n380), .A2(new_n383), .B1(new_n391), .B2(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n393));
  NOR4_X1   g0193(.A1(new_n387), .A2(new_n393), .A3(new_n382), .A4(new_n264), .ZN(new_n394));
  OAI21_X1  g0194(.A(G179), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(G169), .C1(new_n384), .C2(new_n388), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n288), .A2(new_n286), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT68), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(G68), .A3(new_n291), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT73), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n400), .A2(new_n403), .A3(G68), .A4(new_n291), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT74), .B1(new_n287), .B2(G68), .ZN(new_n406));
  XOR2_X1   g0206(.A(new_n406), .B(KEYINPUT12), .Z(new_n407));
  OAI22_X1  g0207(.A1(new_n282), .A2(new_n207), .B1(new_n219), .B2(G68), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n278), .A2(new_n202), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n286), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT11), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n398), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n412), .ZN(new_n414));
  OAI21_X1  g0214(.A(G200), .B1(new_n384), .B2(new_n388), .ZN(new_n415));
  OAI21_X1  g0215(.A(G190), .B1(new_n392), .B2(new_n394), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n400), .A2(G77), .A3(new_n291), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n288), .A2(new_n207), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G20), .A2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT15), .B(G87), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n283), .B2(new_n278), .C1(new_n282), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n286), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n265), .B1(new_n381), .B2(new_n208), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT67), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n254), .A2(G232), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n253), .B(new_n428), .C1(new_n215), .C2(new_n254), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n260), .C1(G107), .C2(new_n253), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n425), .A2(new_n426), .ZN(new_n431));
  INV_X1    g0231(.A(new_n304), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n427), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(KEYINPUT69), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(KEYINPUT69), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n424), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n302), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(G200), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n424), .B(new_n440), .C1(new_n336), .C2(new_n437), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n413), .A2(new_n417), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n370), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G274), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n259), .B(G250), .C1(G1), .C2(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(G116), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n250), .A2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n251), .A2(new_n252), .B1(new_n208), .B2(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n215), .A2(new_n254), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n446), .B(new_n447), .C1(new_n452), .C2(new_n259), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(new_n336), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT19), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n282), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n219), .B1(new_n377), .B2(new_n455), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n209), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n253), .A2(new_n219), .A3(G68), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n460), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n457), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(new_n286), .B1(new_n288), .B2(new_n421), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n218), .A2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n399), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n453), .A2(G200), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n454), .A2(new_n467), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT80), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(G41), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n258), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n445), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n478), .A2(G257), .A3(new_n259), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(new_n254), .C1(new_n319), .C2(new_n320), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT79), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  OAI21_X1  g0282(.A(G250), .B1(new_n319), .B2(new_n320), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G1698), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT79), .B(new_n484), .C1(new_n321), .C2(new_n208), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n482), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n479), .B1(new_n490), .B2(new_n260), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n476), .A2(new_n477), .A3(new_n445), .A4(G274), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(G190), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n287), .A2(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n469), .A2(new_n456), .ZN(new_n495));
  OAI21_X1  g0295(.A(G107), .B1(new_n322), .B2(new_n323), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n456), .A2(new_n459), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n459), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n277), .A2(G77), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n496), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI211_X1 g0305(.A(new_n494), .B(new_n495), .C1(new_n505), .C2(new_n286), .ZN(new_n506));
  INV_X1    g0306(.A(new_n492), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n479), .B(new_n507), .C1(new_n490), .C2(new_n260), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n493), .B(new_n506), .C1(new_n299), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n491), .A2(new_n432), .A3(new_n492), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n494), .B1(new_n505), .B2(new_n286), .ZN(new_n511));
  INV_X1    g0311(.A(new_n495), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n510), .B(new_n513), .C1(G169), .C2(new_n508), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n469), .A2(new_n421), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n467), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n453), .A2(new_n304), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n453), .A2(new_n302), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AND4_X1   g0319(.A1(new_n473), .A2(new_n509), .A3(new_n514), .A4(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n219), .B(G87), .C1(new_n319), .C2(new_n320), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n253), .A2(KEYINPUT85), .A3(new_n219), .A4(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT86), .ZN(new_n526));
  INV_X1    g0326(.A(new_n521), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(KEYINPUT22), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n449), .A2(new_n219), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n219), .A2(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n535), .B(KEYINPUT23), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n530), .A2(new_n534), .A3(new_n531), .A4(new_n536), .ZN(new_n538));
  INV_X1    g0338(.A(new_n533), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n290), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n535), .A2(new_n218), .A3(G13), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT25), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n470), .B2(G107), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n210), .A2(new_n254), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n228), .A2(G1698), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(new_n319), .C2(new_n320), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n260), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n478), .A2(G264), .A3(new_n259), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n492), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n299), .B2(new_n553), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n541), .A2(new_n545), .A3(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n553), .A2(KEYINPUT88), .A3(G169), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT88), .B1(new_n553), .B2(G169), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n551), .A2(G179), .A3(new_n492), .A4(new_n552), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n538), .A2(new_n539), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n538), .A2(new_n539), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n286), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(new_n544), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n489), .B(new_n219), .C1(G33), .C2(new_n456), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n286), .C1(new_n219), .C2(G116), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n399), .A2(KEYINPUT68), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n290), .A2(KEYINPUT68), .A3(new_n287), .ZN(new_n573));
  OAI211_X1 g0373(.A(G116), .B(new_n468), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n287), .A2(G116), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT83), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n254), .A2(G257), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G264), .A2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n319), .C2(new_n320), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n251), .A2(new_n581), .A3(new_n252), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n260), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n478), .A2(G270), .A3(new_n259), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n492), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT82), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT82), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n584), .A3(new_n587), .A4(new_n492), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(G169), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n567), .B1(new_n577), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n585), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G179), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n589), .B2(new_n567), .ZN(new_n595));
  INV_X1    g0395(.A(new_n577), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT84), .B(new_n567), .C1(new_n577), .C2(new_n589), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n586), .A2(new_n588), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G190), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n299), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n596), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n443), .A2(new_n520), .A3(new_n566), .A4(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n358), .A2(new_n359), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n353), .A2(KEYINPUT18), .A3(new_n357), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n439), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n417), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n413), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n608), .B1(new_n613), .B2(new_n352), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n296), .A2(new_n301), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n305), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n514), .A2(new_n509), .A3(new_n473), .ZN(new_n618));
  INV_X1    g0418(.A(new_n555), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n564), .A2(new_n544), .A3(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n620), .C1(new_n565), .C2(new_n599), .ZN(new_n621));
  INV_X1    g0421(.A(new_n519), .ZN(new_n622));
  INV_X1    g0422(.A(new_n514), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n519), .A2(new_n473), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n625), .A3(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n514), .B2(new_n624), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n443), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n617), .A2(new_n631), .ZN(G369));
  NOR2_X1   g0432(.A1(new_n226), .A2(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n218), .ZN(new_n634));
  XNOR2_X1  g0434(.A(KEYINPUT90), .B(KEYINPUT27), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n596), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n604), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n599), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n641), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n640), .B1(new_n541), .B2(new_n545), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n566), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n565), .ZN(new_n649));
  INV_X1    g0449(.A(new_n640), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n620), .B(new_n650), .C1(new_n565), .C2(new_n599), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT91), .Z(G399));
  NOR2_X1   g0455(.A1(new_n460), .A2(G116), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT92), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n227), .A2(G41), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n657), .A2(new_n218), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n223), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT28), .Z(new_n662));
  NAND4_X1  g0462(.A1(new_n566), .A2(new_n520), .A3(new_n604), .A4(new_n650), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n491), .A2(new_n492), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n453), .A2(new_n586), .A3(new_n553), .A4(new_n588), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n432), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT30), .ZN(new_n667));
  AOI211_X1 g0467(.A(new_n479), .B(new_n585), .C1(new_n490), .C2(new_n260), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n559), .A2(new_n453), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n667), .A2(new_n491), .A3(new_n593), .A4(new_n669), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT93), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT93), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n674), .B(new_n666), .C1(new_n670), .C2(new_n671), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n640), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT31), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n663), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n640), .B1(new_n621), .B2(new_n629), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n514), .A2(new_n624), .A3(new_n627), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(KEYINPUT94), .B2(new_n628), .ZN(new_n688));
  AND4_X1   g0488(.A1(KEYINPUT94), .A2(new_n623), .A3(KEYINPUT26), .A4(new_n625), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n519), .B(new_n621), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n686), .B1(new_n690), .B2(new_n650), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n682), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n662), .B1(new_n692), .B2(G1), .ZN(G364));
  AOI21_X1  g0493(.A(new_n218), .B1(new_n633), .B2(G45), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n658), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n646), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(G330), .B2(new_n644), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n224), .B1(G20), .B2(new_n302), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT96), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(G13), .A2(G33), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G20), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n227), .A2(new_n321), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n706), .A2(G355), .B1(new_n448), .B2(new_n227), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT95), .Z(new_n708));
  NAND2_X1  g0508(.A1(new_n660), .A2(new_n444), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n244), .B2(new_n444), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n227), .A2(new_n253), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n705), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n696), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n219), .A2(G190), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n299), .A2(G179), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT99), .Z(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n459), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G159), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT32), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n321), .B1(new_n724), .B2(KEYINPUT32), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n219), .A2(new_n336), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n717), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G87), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n336), .A2(G179), .A3(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n219), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G97), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n725), .A2(new_n726), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n716), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n432), .A2(G200), .A3(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n720), .B(new_n735), .C1(G77), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n304), .A2(G200), .A3(new_n727), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT98), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n739), .A2(KEYINPUT98), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n304), .A2(new_n299), .A3(new_n727), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT97), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G50), .A2(new_n744), .B1(new_n751), .B2(G58), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n432), .A2(new_n299), .A3(new_n736), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n738), .B(new_n752), .C1(new_n214), .C2(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT100), .B(G326), .Z(new_n756));
  AOI22_X1  g0556(.A1(G322), .A2(new_n751), .B1(new_n744), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n321), .B1(new_n728), .B2(new_n581), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT101), .ZN(new_n759));
  INV_X1    g0559(.A(new_n737), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(KEYINPUT101), .B2(new_n758), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(new_n753), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n723), .A2(G329), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n719), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G294), .B2(new_n733), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n757), .A2(new_n759), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n715), .B1(new_n770), .B2(new_n701), .ZN(new_n771));
  INV_X1    g0571(.A(new_n704), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n714), .B(new_n771), .C1(new_n644), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n698), .A2(new_n773), .ZN(G396));
  INV_X1    g0574(.A(KEYINPUT104), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n609), .A2(KEYINPUT103), .A3(new_n640), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n439), .B(new_n441), .C1(new_n424), .C2(new_n650), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT103), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n439), .B2(new_n650), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n684), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n683), .A2(new_n780), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n775), .B1(new_n785), .B2(new_n682), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n682), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(KEYINPUT104), .A3(new_n681), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n786), .A2(new_n715), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n719), .A2(new_n214), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n253), .B1(new_n728), .B2(new_n202), .C1(new_n732), .C2(new_n313), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n744), .A2(G137), .B1(G159), .B2(new_n737), .ZN(new_n792));
  INV_X1    g0592(.A(G143), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(new_n276), .B2(new_n754), .C1(new_n793), .C2(new_n750), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT34), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n790), .B(new_n791), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n723), .A2(G132), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n795), .C2(new_n794), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n719), .A2(new_n209), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G311), .B2(new_n723), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT102), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n734), .B1(new_n766), .B2(new_n754), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n321), .B1(new_n459), .B2(new_n728), .C1(new_n760), .C2(new_n448), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n800), .A2(new_n801), .B1(G294), .B2(new_n751), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(new_n581), .C2(new_n743), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n715), .B1(new_n807), .B2(new_n701), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n701), .A2(new_n702), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(G77), .B2(new_n810), .C1(new_n703), .C2(new_n780), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n789), .A2(new_n811), .ZN(G384));
  NAND4_X1  g0612(.A1(new_n673), .A2(KEYINPUT31), .A3(new_n640), .A4(new_n675), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n663), .A2(new_n678), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n412), .A2(new_n640), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n413), .A2(new_n417), .A3(new_n815), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n412), .B(new_n640), .C1(new_n817), .C2(new_n398), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n814), .A2(new_n819), .A3(new_n780), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT108), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n349), .A2(new_n350), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n349), .A2(new_n350), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n348), .A2(KEYINPUT108), .A3(new_n351), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n608), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n638), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n353), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n358), .A2(new_n829), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n347), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n327), .A2(new_n340), .A3(new_n346), .ZN(new_n835));
  INV_X1    g0635(.A(new_n832), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n358), .A2(new_n829), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT38), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n342), .A2(new_n343), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n327), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n828), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n607), .A2(KEYINPUT76), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n358), .A2(KEYINPUT77), .A3(new_n359), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n362), .B1(new_n361), .B2(KEYINPUT18), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n361), .A2(new_n365), .A3(KEYINPUT18), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n823), .A2(new_n824), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n841), .B1(new_n357), .B2(new_n828), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n835), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n837), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT110), .B1(new_n839), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT38), .B(new_n853), .C1(new_n369), .C2(new_n842), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT110), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n827), .A2(new_n830), .B1(new_n837), .B2(new_n834), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(KEYINPUT38), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n821), .A2(new_n857), .A3(KEYINPUT40), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n855), .B1(new_n849), .B2(new_n854), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n820), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n443), .A2(new_n814), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n868), .B(new_n869), .Z(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(G330), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n443), .B1(new_n685), .B2(new_n691), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n617), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT109), .Z(new_n874));
  XNOR2_X1  g0674(.A(new_n871), .B(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n439), .A2(new_n640), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n683), .B2(new_n780), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n858), .A2(new_n864), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n819), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n606), .A2(new_n607), .A3(new_n638), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n398), .A2(new_n412), .A3(new_n650), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT107), .Z(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n839), .B2(new_n856), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n858), .A2(new_n864), .A3(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n880), .B(new_n881), .C1(new_n883), .C2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n875), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n875), .A2(new_n888), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n889), .B(new_n890), .C1(new_n218), .C2(new_n633), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n448), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n224), .A2(new_n219), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n892), .B(new_n893), .C1(KEYINPUT35), .C2(new_n502), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI21_X1  g0695(.A(G77), .B1(new_n313), .B2(new_n214), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n896), .A2(new_n223), .B1(G50), .B2(new_n214), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G1), .A3(new_n226), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT105), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n891), .A2(new_n895), .A3(new_n899), .ZN(G367));
  NAND2_X1  g0700(.A1(new_n509), .A2(new_n514), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n506), .B2(new_n650), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n514), .B2(new_n650), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(new_n653), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT45), .Z(new_n906));
  INV_X1    g0706(.A(new_n652), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n653), .A2(new_n902), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT44), .Z(new_n909));
  OR3_X1    g0709(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n906), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n643), .A2(new_n640), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n566), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n651), .B2(new_n913), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(new_n645), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n692), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n658), .B(KEYINPUT41), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n695), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n650), .B1(new_n467), .B2(new_n471), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n622), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n624), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT112), .Z(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(KEYINPUT113), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n925));
  OR3_X1    g0725(.A1(new_n914), .A2(KEYINPUT42), .A3(new_n903), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n514), .B1(new_n903), .B2(new_n649), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n650), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT42), .B1(new_n914), .B2(new_n903), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n924), .A2(KEYINPUT113), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n931), .A2(new_n933), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n907), .A2(new_n904), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n937), .B(new_n938), .Z(new_n939));
  OR2_X1    g0739(.A1(new_n919), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n728), .A2(new_n448), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT46), .ZN(new_n942));
  INV_X1    g0742(.A(new_n718), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n253), .B1(new_n943), .B2(G97), .ZN(new_n944));
  INV_X1    g0744(.A(G294), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n944), .B1(new_n754), .B2(new_n945), .C1(new_n766), .C2(new_n760), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n942), .B(new_n946), .C1(G107), .C2(new_n733), .ZN(new_n947));
  XOR2_X1   g0747(.A(KEYINPUT114), .B(G311), .Z(new_n948));
  AOI22_X1  g0748(.A1(G303), .A2(new_n751), .B1(new_n744), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(G317), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n947), .B(new_n949), .C1(new_n950), .C2(new_n722), .ZN(new_n951));
  INV_X1    g0751(.A(G159), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n202), .A2(new_n760), .B1(new_n754), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G58), .A2(new_n729), .B1(new_n723), .B2(G137), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(KEYINPUT115), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n253), .B1(new_n718), .B2(new_n207), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n732), .A2(new_n214), .ZN(new_n957));
  NOR4_X1   g0757(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G143), .A2(new_n744), .B1(new_n751), .B2(G150), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n954), .A2(KEYINPUT115), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n951), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT47), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n715), .B1(new_n963), .B2(new_n701), .ZN(new_n964));
  INV_X1    g0764(.A(new_n227), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n705), .B1(new_n965), .B2(new_n421), .C1(new_n240), .C2(new_n712), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(new_n772), .C2(new_n922), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n940), .A2(new_n967), .ZN(G387));
  AOI21_X1  g0768(.A(new_n712), .B1(new_n236), .B2(G45), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n657), .B2(new_n706), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n444), .A3(new_n972), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n657), .B(new_n973), .C1(G68), .C2(G77), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n970), .A2(new_n974), .B1(G107), .B2(new_n965), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n715), .B1(new_n975), .B2(new_n705), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT116), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n723), .A2(new_n756), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n751), .A2(G317), .B1(G303), .B2(new_n737), .ZN(new_n979));
  INV_X1    g0779(.A(G322), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n743), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n753), .B2(new_n948), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT48), .Z(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n766), .B2(new_n732), .C1(new_n945), .C2(new_n728), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT49), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n253), .B(new_n978), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n985), .B2(new_n984), .C1(new_n448), .C2(new_n718), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G50), .A2(new_n751), .B1(new_n744), .B2(G159), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n214), .A2(new_n760), .B1(new_n754), .B2(new_n283), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n253), .B1(new_n728), .B2(new_n207), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT117), .B(G150), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n723), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n421), .B2(new_n732), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n988), .B(new_n994), .C1(new_n456), .C2(new_n719), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n977), .B1(new_n651), .B2(new_n772), .C1(new_n996), .C2(new_n700), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n916), .A2(new_n694), .ZN(new_n998));
  INV_X1    g0798(.A(new_n692), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(new_n916), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n916), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n658), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n998), .A3(new_n1002), .ZN(G393));
  OAI22_X1  g0803(.A1(new_n276), .A2(new_n743), .B1(new_n750), .B2(new_n952), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT51), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n321), .B1(new_n729), .B2(G68), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n733), .A2(G77), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n793), .C2(new_n722), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1008), .B(new_n799), .C1(new_n341), .C2(new_n737), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1005), .B(new_n1009), .C1(new_n202), .C2(new_n754), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n761), .A2(new_n750), .B1(new_n743), .B2(new_n950), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT52), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n253), .B1(new_n729), .B2(G283), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n448), .B2(new_n732), .C1(new_n980), .C2(new_n722), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n720), .B(new_n1014), .C1(G294), .C2(new_n737), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1012), .B(new_n1015), .C1(new_n581), .C2(new_n754), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n715), .B1(new_n1017), .B2(new_n701), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n705), .B1(new_n456), .B2(new_n965), .C1(new_n247), .C2(new_n712), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n772), .C2(new_n904), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n912), .B2(new_n694), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n912), .A2(new_n1000), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n658), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n912), .B2(new_n1000), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(G390));
  NAND3_X1  g0826(.A1(new_n443), .A2(G330), .A3(new_n814), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n616), .A2(new_n305), .A3(new_n872), .A4(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n690), .A2(new_n650), .A3(new_n780), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n876), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n682), .A2(new_n780), .A3(new_n819), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n814), .A2(KEYINPUT119), .A3(G330), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT119), .B1(new_n814), .B2(G330), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n781), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1031), .B(new_n1032), .C1(new_n1035), .C2(new_n819), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n821), .A2(G330), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n819), .B1(new_n682), .B2(new_n780), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n878), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1028), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n819), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n883), .B1(new_n877), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n887), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n857), .A2(new_n861), .A3(new_n883), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1041), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1037), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1043), .B(new_n1032), .C1(new_n1046), .C2(new_n1045), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT118), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1052), .A2(KEYINPUT118), .A3(new_n1043), .A4(new_n1032), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1040), .A2(new_n1048), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(new_n658), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1058), .B2(new_n1028), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1056), .A2(new_n694), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n887), .A2(new_n702), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n253), .B1(new_n723), .B2(G294), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1007), .A2(new_n1063), .A3(new_n730), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1064), .B(new_n790), .C1(G97), .C2(new_n737), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G116), .A2(new_n751), .B1(new_n744), .B2(G283), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n459), .C2(new_n754), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G128), .A2(new_n744), .B1(new_n751), .B2(G132), .ZN(new_n1068));
  INV_X1    g0868(.A(G125), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n253), .B1(new_n722), .B2(new_n1069), .C1(new_n202), .C2(new_n718), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT120), .ZN(new_n1071));
  INV_X1    g0871(.A(G137), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n754), .A2(new_n1072), .B1(new_n952), .B2(new_n732), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT54), .B(G143), .Z(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n737), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1068), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n729), .A2(new_n991), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1067), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n715), .B1(new_n1079), .B2(new_n701), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1062), .B(new_n1080), .C1(new_n341), .C2(new_n810), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1061), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1060), .A2(new_n1083), .ZN(G378));
  INV_X1    g0884(.A(KEYINPUT124), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT123), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n857), .A2(new_n861), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n814), .A2(new_n819), .A3(KEYINPUT40), .A4(new_n780), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n866), .B(G330), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT55), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n306), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n296), .A2(new_n301), .A3(new_n305), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT55), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n293), .A2(new_n828), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT56), .Z(new_n1095));
  AND3_X1   g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1089), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n862), .A2(new_n1098), .A3(G330), .A4(new_n866), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n888), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1086), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(KEYINPUT123), .B(new_n888), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1100), .A2(new_n888), .A3(new_n1101), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT122), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT122), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1100), .A2(new_n1109), .A3(new_n888), .A4(new_n1101), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT57), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1028), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1107), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1023), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1098), .A2(new_n702), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n809), .A2(new_n202), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n753), .A2(G132), .B1(new_n729), .B2(new_n1074), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1072), .B2(new_n760), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G128), .B2(new_n751), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n1069), .B2(new_n743), .C1(new_n276), .C2(new_n732), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n250), .B1(new_n718), .B2(new_n952), .ZN(new_n1129));
  AOI211_X1 g0929(.A(G41), .B(new_n1129), .C1(G124), .C2(new_n723), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n202), .B1(new_n319), .B2(G41), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n321), .B1(new_n754), .B2(new_n456), .C1(new_n421), .C2(new_n760), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G116), .B2(new_n744), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G58), .A2(new_n943), .B1(new_n723), .B2(G283), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n207), .B2(new_n728), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1139), .A2(G41), .A3(new_n957), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(new_n459), .C2(new_n750), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT58), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1134), .A2(new_n1135), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n715), .B1(new_n1143), .B2(new_n701), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1122), .A2(new_n1123), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1117), .A2(KEYINPUT123), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1102), .A2(new_n1086), .A3(new_n1103), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1111), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1149), .B2(new_n695), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1085), .B1(new_n1121), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1119), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1153));
  OAI211_X1 g0953(.A(KEYINPUT124), .B(new_n1150), .C1(new_n1153), .C2(new_n1023), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(G375));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n253), .B1(new_n722), .B2(new_n1157), .C1(new_n313), .C2(new_n718), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n732), .A2(new_n202), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n753), .A2(new_n1074), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n760), .B2(new_n276), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G132), .C2(new_n744), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n1072), .B2(new_n750), .C1(new_n952), .C2(new_n728), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n754), .A2(new_n448), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n760), .A2(new_n459), .B1(new_n719), .B2(new_n207), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n321), .B1(new_n722), .B2(new_n581), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n732), .A2(new_n421), .B1(new_n728), .B2(new_n456), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n766), .B2(new_n750), .C1(new_n945), .C2(new_n743), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1164), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n715), .B1(new_n1171), .B2(new_n701), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n819), .B2(new_n703), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n214), .B2(new_n809), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n694), .B(KEYINPUT125), .Z(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1057), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1028), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n918), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1178), .B2(new_n1040), .ZN(G381));
  OAI211_X1 g0979(.A(new_n1025), .B(new_n967), .C1(new_n919), .C2(new_n939), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1082), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1152), .A2(new_n1181), .A3(new_n1154), .ZN(new_n1182));
  INV_X1    g0982(.A(G396), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n997), .A2(new_n1183), .A3(new_n998), .A4(new_n1002), .ZN(new_n1184));
  OR2_X1    g0984(.A1(G381), .A2(G384), .ZN(new_n1185));
  OR4_X1    g0985(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .A4(new_n1185), .ZN(G407));
  OAI211_X1 g0986(.A(G407), .B(G213), .C1(G343), .C2(new_n1182), .ZN(G409));
  AOI21_X1  g0987(.A(new_n1025), .B1(new_n940), .B2(new_n967), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(G393), .A2(G396), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1184), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1191), .A3(new_n1180), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1180), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1184), .B(new_n1190), .C1(new_n1188), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G378), .B(new_n1150), .C1(new_n1153), .C2(new_n1023), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1118), .A2(new_n1175), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1145), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1106), .A2(new_n1111), .B1(new_n1113), .B2(new_n1054), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(new_n918), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n1201), .B2(G378), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1149), .A2(new_n918), .A3(new_n1114), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n1145), .A3(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(KEYINPUT126), .A3(new_n1181), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1196), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n639), .A2(G213), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT60), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1177), .B1(new_n1040), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT127), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1177), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1023), .B1(new_n1213), .B2(KEYINPUT60), .ZN(new_n1214));
  OAI211_X1 g1014(.A(KEYINPUT127), .B(new_n1177), .C1(new_n1040), .C2(new_n1209), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G384), .B1(new_n1216), .B2(new_n1176), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(G384), .A3(new_n1176), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n639), .A2(G213), .A3(G2897), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1220), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1216), .A2(G384), .A3(new_n1176), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n1217), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1208), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1223), .A2(new_n1217), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1206), .A2(new_n1228), .A3(new_n1207), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT62), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT62), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT61), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1195), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1229), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1225), .B1(new_n1207), .B2(new_n1206), .ZN(new_n1236));
  OAI21_X1  g1036(.A(KEYINPUT63), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT63), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1195), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1232), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1240), .ZN(G405));
  OAI21_X1  g1041(.A(G378), .B1(new_n1121), .B2(new_n1151), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1195), .A2(new_n1182), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1195), .B1(new_n1182), .B2(new_n1242), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1228), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1182), .A2(new_n1242), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1194), .A3(new_n1192), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1228), .B1(new_n1249), .B2(new_n1243), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1247), .A2(new_n1250), .ZN(G402));
endmodule


