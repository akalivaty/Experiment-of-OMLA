//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT25), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT23), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT65), .B(G169gat), .Z(new_n225));
  NAND4_X1  g024(.A1(new_n225), .A2(KEYINPUT66), .A3(KEYINPUT23), .A4(new_n214), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n213), .A2(new_n220), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n228));
  OR2_X1    g027(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n229), .A2(KEYINPUT27), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT27), .B(G183gat), .Z(new_n234));
  OAI21_X1  g033(.A(KEYINPUT28), .B1(new_n234), .B2(G190gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n212), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(new_n203), .A3(new_n235), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n242));
  AOI21_X1  g041(.A(G190gat), .B1(new_n229), .B2(new_n230), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n205), .A2(new_n206), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n212), .B(new_n242), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n222), .B(KEYINPUT67), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT25), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n241), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G226gat), .ZN(new_n249));
  INV_X1    g048(.A(G233gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(KEYINPUT29), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n251), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n227), .A2(new_n241), .A3(new_n247), .A4(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n258), .A3(new_n262), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n266), .A2(KEYINPUT73), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT73), .B1(new_n266), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n202), .B1(new_n257), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n256), .ZN(new_n274));
  INV_X1    g073(.A(new_n270), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n271), .A2(new_n273), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT74), .B1(new_n274), .B2(new_n275), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n202), .B(new_n270), .C1(new_n254), .C2(new_n256), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n286), .A2(KEYINPUT75), .A3(new_n273), .A4(new_n280), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT76), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n281), .A2(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n273), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n279), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n283), .A2(new_n287), .A3(new_n294), .A4(new_n288), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT69), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n301), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n303), .B(new_n304), .C1(KEYINPUT1), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(G120gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(G113gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n314), .A2(KEYINPUT70), .A3(new_n304), .A4(new_n303), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n302), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G148gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G141gat), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT2), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n326), .B1(new_n325), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n318), .B1(new_n308), .B2(new_n315), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n298), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n330), .B2(new_n331), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n329), .ZN(new_n342));
  INV_X1    g141(.A(new_n326), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT4), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n339), .B1(new_n349), .B2(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT71), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n353), .B(new_n318), .C1(new_n308), .C2(new_n315), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT4), .B(new_n332), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n350), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n340), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  NOR2_X1   g162(.A1(new_n335), .A2(new_n348), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n336), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n332), .B1(new_n352), .B2(new_n354), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n364), .B(new_n366), .C1(new_n367), .C2(new_n365), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n297), .A2(new_n339), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n358), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n363), .B1(new_n358), .B2(new_n370), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(KEYINPUT6), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n296), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT81), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(new_n373), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT80), .ZN(new_n383));
  INV_X1    g182(.A(new_n376), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n378), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n296), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n272), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n332), .B1(new_n392), .B2(new_n345), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n272), .B1(new_n347), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n270), .B1(new_n391), .B2(new_n347), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n396), .A2(new_n393), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n399));
  AND2_X1   g198(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  INV_X1    g201(.A(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n398), .A2(G22gat), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(KEYINPUT84), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n398), .B(G22gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n320), .A2(new_n353), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n227), .A2(new_n241), .A3(new_n247), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n248), .B1(new_n352), .B2(new_n354), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT64), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT34), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT72), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n419), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(KEYINPUT34), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n416), .A2(new_n417), .B1(G227gat), .B2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n427), .A2(KEYINPUT72), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n423), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT32), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n424), .A3(KEYINPUT34), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT72), .B1(new_n427), .B2(new_n428), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n432), .A3(new_n423), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n434), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n423), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n447), .B(new_n433), .C1(new_n442), .C2(new_n443), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n432), .B1(new_n444), .B2(new_n423), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n440), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n412), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n381), .A2(new_n389), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT87), .B1(new_n382), .B2(new_n376), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n384), .A2(new_n455), .A3(new_n373), .A4(new_n371), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(new_n378), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(new_n296), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n451), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n409), .A2(new_n411), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n462));
  AOI211_X1 g261(.A(KEYINPUT81), .B(new_n462), .C1(new_n378), .C2(new_n386), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n388), .B1(new_n387), .B2(new_n296), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n450), .A2(KEYINPUT36), .A3(new_n446), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT36), .B1(new_n450), .B2(new_n446), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  INV_X1    g268(.A(new_n364), .ZN(new_n470));
  INV_X1    g269(.A(new_n366), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n333), .B1(new_n413), .B2(new_n415), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(KEYINPUT4), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n473), .A2(new_n474), .A3(new_n339), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n473), .B2(new_n339), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT85), .B1(new_n368), .B2(new_n338), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n474), .A3(new_n339), .ZN(new_n479));
  INV_X1    g278(.A(new_n337), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n469), .B1(new_n480), .B2(new_n338), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n482), .A3(new_n363), .ZN(new_n483));
  NOR2_X1   g282(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n482), .A3(new_n363), .A4(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(new_n384), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n461), .B1(new_n488), .B2(new_n462), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n454), .A2(new_n456), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n286), .A2(new_n491), .A3(new_n273), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n274), .A2(new_n272), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(KEYINPUT37), .C1(new_n274), .C2(new_n270), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n279), .A4(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT88), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n292), .A2(KEYINPUT37), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n279), .A3(new_n492), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT38), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n501), .A2(new_n283), .A3(new_n287), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n490), .A2(new_n498), .A3(new_n502), .A4(new_n378), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n468), .B1(new_n489), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n453), .A2(new_n460), .B1(new_n465), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G15gat), .B(G22gat), .Z(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  OR3_X1    g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n510), .C1(KEYINPUT16), .C2(new_n506), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(G8gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(G8gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT89), .ZN(new_n520));
  OR3_X1    g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(KEYINPUT90), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n522), .B2(KEYINPUT90), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n518), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n521), .B(KEYINPUT91), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n520), .ZN(new_n531));
  INV_X1    g330(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n527), .A4(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n529), .A2(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT17), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n514), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n514), .A2(new_n538), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR4_X1   g344(.A1(new_n540), .A2(new_n541), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n514), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n535), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n542), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n544), .B(KEYINPUT13), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT94), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n539), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n547), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n544), .A3(new_n542), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n555), .B(new_n552), .C1(new_n558), .C2(new_n541), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n540), .A2(new_n545), .A3(new_n543), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT93), .B1(new_n560), .B2(KEYINPUT18), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n562), .A3(new_n541), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n554), .A2(new_n559), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G113gat), .B(G141gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT11), .B(G169gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT12), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n546), .A2(new_n553), .A3(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(KEYINPUT18), .B2(new_n560), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n571), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT96), .B1(new_n505), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n465), .A2(new_n504), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n452), .A2(KEYINPUT35), .B1(new_n451), .B2(new_n459), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n580), .B(new_n577), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  XNOR2_X1  g387(.A(G57gat), .B(G64gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n547), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(new_n207), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(KEYINPUT21), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n595), .B(G183gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G211gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n599), .A2(new_n601), .A3(G231gat), .A4(G233gat), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n604), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n587), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n608), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n606), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n586), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G99gat), .B(G106gat), .Z(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n617), .A2(KEYINPUT98), .B1(KEYINPUT8), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(G85gat), .A3(G92gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT7), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n619), .B(new_n622), .C1(G85gat), .C2(G92gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n537), .B2(new_n539), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n628), .A2(KEYINPUT99), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(KEYINPUT99), .B2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n538), .A2(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G190gat), .B(G218gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n630), .A2(new_n629), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n642), .A3(new_n637), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n616), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n625), .A2(new_n626), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n594), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n627), .A2(new_n593), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(KEYINPUT101), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT101), .B1(new_n627), .B2(new_n593), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(KEYINPUT10), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G230gat), .ZN(new_n658));
  OAI22_X1  g457(.A1(new_n655), .A2(new_n657), .B1(new_n658), .B2(new_n250), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n653), .B(new_n650), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n250), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n647), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n647), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n585), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n387), .B(KEYINPUT103), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT104), .B(G1gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1324gat));
  NOR2_X1   g481(.A1(new_n676), .A2(new_n296), .ZN(new_n683));
  NAND2_X1  g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  OR2_X1    g483(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  INV_X1    g488(.A(G8gat), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n688), .B(new_n689), .C1(new_n690), .C2(new_n683), .ZN(G1325gat));
  AND3_X1   g490(.A1(new_n677), .A2(G15gat), .A3(new_n468), .ZN(new_n692));
  INV_X1    g491(.A(new_n446), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n441), .B1(new_n434), .B2(new_n445), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(G15gat), .B1(new_n677), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n692), .A2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n461), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n616), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n669), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n585), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(new_n524), .A3(new_n646), .A4(new_n679), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n571), .A2(new_n574), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  INV_X1    g506(.A(new_n645), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n642), .B1(new_n636), .B2(new_n637), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n453), .A2(new_n460), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n581), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n505), .C2(new_n710), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n646), .A2(new_n713), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n412), .B1(new_n381), .B2(new_n389), .ZN(new_n720));
  INV_X1    g519(.A(new_n467), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n450), .A2(new_n446), .A3(KEYINPUT36), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n501), .A2(new_n283), .A3(new_n287), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n457), .A2(new_n724), .A3(new_n497), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n485), .A2(new_n384), .A3(new_n487), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n412), .B1(new_n726), .B2(new_n296), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n723), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n719), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n465), .A2(new_n504), .A3(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n718), .B1(new_n731), .B2(new_n583), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n711), .A2(new_n729), .A3(KEYINPUT107), .A4(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n717), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n706), .B(new_n702), .C1(new_n716), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G29gat), .B1(new_n735), .B2(new_n678), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n705), .A2(new_n736), .ZN(G1328gat));
  AND2_X1   g536(.A1(new_n703), .A2(new_n646), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n525), .A3(new_n462), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  OAI21_X1  g539(.A(G36gat), .B1(new_n735), .B2(new_n296), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n738), .A2(new_n742), .A3(new_n525), .A4(new_n462), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(G1329gat));
  NAND4_X1  g543(.A1(new_n585), .A2(new_n695), .A3(new_n646), .A4(new_n702), .ZN(new_n745));
  INV_X1    g544(.A(G43gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n468), .A2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n735), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT48), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n585), .A2(new_n461), .A3(new_n646), .A4(new_n702), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n403), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n461), .A2(G50gat), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n752), .B(new_n754), .C1(new_n735), .C2(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n751), .A2(KEYINPUT48), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1331gat));
  INV_X1    g557(.A(new_n706), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n647), .A2(new_n759), .A3(new_n669), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n732), .B2(new_n733), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n679), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n462), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n765), .B(new_n766), .Z(G1333gat));
  NAND2_X1  g566(.A1(new_n761), .A2(new_n695), .ZN(new_n768));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n723), .A2(new_n769), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n761), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n761), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n775), .B(new_n776), .Z(G1334gat));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n461), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT111), .B(G78gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n701), .A2(new_n706), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n646), .B(new_n781), .C1(new_n731), .C2(new_n583), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT51), .ZN(new_n783));
  OR4_X1    g582(.A1(G85gat), .A2(new_n783), .A3(new_n670), .A4(new_n678), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n669), .B(new_n781), .C1(new_n716), .C2(new_n734), .ZN(new_n785));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n678), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1336gat));
  OAI21_X1  g586(.A(G92gat), .B1(new_n785), .B2(new_n296), .ZN(new_n788));
  INV_X1    g587(.A(new_n783), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n670), .A2(G92gat), .A3(new_n296), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT112), .Z(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n788), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1337gat));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n785), .A2(new_n798), .A3(new_n723), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n785), .B2(new_n723), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(G99gat), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(G99gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n695), .A2(new_n802), .A3(new_n669), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT114), .Z(new_n804));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(G1338gat));
  OAI21_X1  g605(.A(G106gat), .B1(new_n785), .B2(new_n412), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n412), .A2(G106gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n669), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1339gat));
  INV_X1    g613(.A(new_n568), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n544), .B1(new_n557), .B2(new_n542), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n549), .A2(new_n551), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n574), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n669), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n661), .B(new_n656), .C1(new_n660), .C2(KEYINPUT10), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n659), .A2(new_n821), .A3(KEYINPUT54), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  OAI221_X1 g622(.A(new_n823), .B1(new_n658), .B2(new_n250), .C1(new_n655), .C2(new_n657), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n666), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n666), .A4(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n667), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n820), .B1(new_n759), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n710), .ZN(new_n831));
  INV_X1    g630(.A(new_n829), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n646), .A2(new_n819), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n701), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n616), .A2(new_n646), .A3(new_n706), .A4(new_n669), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n679), .A2(new_n296), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n451), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n578), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n706), .A2(new_n310), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(G1340gat));
  NOR2_X1   g641(.A1(new_n839), .A2(new_n670), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(new_n312), .ZN(G1341gat));
  NOR2_X1   g643(.A1(new_n839), .A2(new_n616), .ZN(new_n845));
  XOR2_X1   g644(.A(KEYINPUT115), .B(G127gat), .Z(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(G1342gat));
  AOI21_X1  g646(.A(new_n839), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n646), .ZN(new_n849));
  NOR2_X1   g648(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT116), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n849), .B(new_n851), .ZN(G1343gat));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n825), .A2(new_n853), .A3(new_n826), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n825), .B2(new_n826), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n828), .A2(new_n667), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n577), .A2(new_n858), .B1(new_n669), .B2(new_n819), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n833), .B1(new_n859), .B2(new_n646), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n835), .B1(new_n860), .B2(new_n616), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n412), .ZN(new_n862));
  INV_X1    g661(.A(new_n837), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n723), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n834), .A2(new_n835), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n461), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n862), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n323), .B1(new_n870), .B2(new_n706), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n468), .A2(new_n412), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n866), .A2(new_n863), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(G141gat), .A3(new_n578), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT58), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n577), .A3(new_n868), .A4(new_n865), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(G141gat), .B2(new_n878), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n880));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(G141gat), .ZN(new_n882));
  INV_X1    g681(.A(new_n876), .ZN(new_n883));
  AND4_X1   g682(.A1(KEYINPUT120), .A2(new_n882), .A3(new_n883), .A4(new_n880), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n877), .B1(new_n881), .B2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(new_n875), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n321), .A3(new_n669), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n706), .A2(KEYINPUT95), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n856), .A2(new_n857), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n854), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n646), .B1(new_n893), .B2(new_n820), .ZN(new_n894));
  INV_X1    g693(.A(new_n833), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT122), .B(new_n833), .C1(new_n859), .C2(new_n646), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n616), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n672), .A2(new_n578), .A3(new_n674), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n461), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n461), .C1(new_n834), .C2(new_n835), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT121), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n669), .B(new_n865), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n888), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n321), .C1(new_n870), .C2(new_n669), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n887), .B1(new_n905), .B2(new_n906), .ZN(G1345gat));
  AOI21_X1  g706(.A(G155gat), .B1(new_n886), .B2(new_n701), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n616), .A2(new_n327), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n870), .B2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(new_n328), .B1(new_n875), .B2(new_n710), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n646), .A2(G162gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n869), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT123), .Z(G1347gat));
  NAND2_X1  g713(.A1(new_n451), .A2(new_n462), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n866), .A2(new_n916), .A3(new_n678), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n836), .B2(new_n679), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n225), .A3(new_n706), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n451), .A2(new_n462), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n866), .A2(new_n678), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n578), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(G1348gat));
  NOR3_X1   g723(.A1(new_n922), .A2(new_n214), .A3(new_n670), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n919), .A2(new_n669), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n214), .ZN(G1349gat));
  NOR2_X1   g726(.A1(new_n616), .A2(new_n234), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n919), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n229), .B(new_n230), .C1(new_n922), .C2(new_n616), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n919), .A2(new_n208), .A3(new_n646), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n922), .B2(new_n710), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  OR2_X1    g737(.A1(new_n901), .A2(new_n903), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n678), .A2(new_n462), .A3(new_n723), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT126), .Z(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n577), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G197gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n872), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n917), .B2(new_n918), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n462), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n759), .A2(G197gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n945), .A2(new_n949), .A3(new_n462), .A4(new_n669), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n939), .A2(new_n669), .A3(new_n941), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n951), .B(new_n952), .C1(new_n953), .C2(new_n949), .ZN(G1353gat));
  NAND4_X1  g753(.A1(new_n945), .A2(new_n260), .A3(new_n462), .A4(new_n701), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n701), .B(new_n941), .C1(new_n901), .C2(new_n903), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  AND3_X1   g758(.A1(new_n939), .A2(new_n646), .A3(new_n941), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n646), .A2(new_n261), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n960), .A2(new_n261), .B1(new_n946), .B2(new_n961), .ZN(G1355gat));
endmodule


