

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759;

  OR2_X1 U374 ( .A1(n392), .A2(n390), .ZN(n514) );
  NOR2_X1 U375 ( .A1(n565), .A2(n566), .ZN(n665) );
  XNOR2_X1 U376 ( .A(n453), .B(KEYINPUT45), .ZN(n673) );
  XNOR2_X1 U377 ( .A(n381), .B(n360), .ZN(n553) );
  BUF_X1 U378 ( .A(n745), .Z(n425) );
  XOR2_X1 U379 ( .A(n427), .B(KEYINPUT30), .Z(n352) );
  AND2_X4 U380 ( .A1(n638), .A2(n639), .ZN(n725) );
  XNOR2_X2 U381 ( .A(n520), .B(G134), .ZN(n529) );
  OR2_X2 U382 ( .A1(n710), .A2(n611), .ZN(n379) );
  INV_X2 U383 ( .A(n692), .ZN(n383) );
  NOR2_X1 U384 ( .A1(n707), .A2(G953), .ZN(n502) );
  NAND2_X1 U385 ( .A1(n479), .A2(n423), .ZN(n478) );
  XNOR2_X1 U386 ( .A(n480), .B(n364), .ZN(n479) );
  AND2_X1 U387 ( .A1(n673), .A2(n477), .ZN(n461) );
  XNOR2_X1 U388 ( .A(n564), .B(n428), .ZN(n759) );
  NOR2_X1 U389 ( .A1(n563), .A2(n588), .ZN(n564) );
  INV_X1 U390 ( .A(n695), .ZN(n612) );
  XNOR2_X1 U391 ( .A(n610), .B(n579), .ZN(n689) );
  OR2_X1 U392 ( .A1(n642), .A2(G902), .ZN(n381) );
  XNOR2_X1 U393 ( .A(n742), .B(G146), .ZN(n507) );
  XNOR2_X1 U394 ( .A(n529), .B(n488), .ZN(n742) );
  XNOR2_X1 U395 ( .A(KEYINPUT0), .B(KEYINPUT68), .ZN(n595) );
  INV_X1 U396 ( .A(KEYINPUT40), .ZN(n428) );
  XOR2_X1 U397 ( .A(G125), .B(G146), .Z(n521) );
  INV_X1 U398 ( .A(KEYINPUT69), .ZN(n415) );
  INV_X2 U399 ( .A(G953), .ZN(n745) );
  XNOR2_X1 U400 ( .A(n598), .B(n476), .ZN(n405) );
  XNOR2_X1 U401 ( .A(n416), .B(n517), .ZN(n519) );
  XNOR2_X2 U402 ( .A(n513), .B(n512), .ZN(n610) );
  NAND2_X1 U403 ( .A1(n439), .A2(n437), .ZN(n376) );
  XNOR2_X1 U404 ( .A(n438), .B(KEYINPUT77), .ZN(n437) );
  AND2_X1 U405 ( .A1(n575), .A2(n440), .ZN(n439) );
  NAND2_X1 U406 ( .A1(n448), .A2(n445), .ZN(n444) );
  XNOR2_X1 U407 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n497) );
  INV_X1 U408 ( .A(KEYINPUT85), .ZN(n634) );
  NAND2_X1 U409 ( .A1(n420), .A2(n633), .ZN(n453) );
  XNOR2_X1 U410 ( .A(n455), .B(n454), .ZN(n420) );
  OR2_X1 U411 ( .A1(n505), .A2(G902), .ZN(n370) );
  AND2_X1 U412 ( .A1(n466), .A2(n464), .ZN(n426) );
  AND2_X1 U413 ( .A1(n559), .A2(n528), .ZN(n465) );
  XNOR2_X1 U414 ( .A(G113), .B(G131), .ZN(n540) );
  NAND2_X1 U415 ( .A1(n745), .A2(G224), .ZN(n416) );
  NOR2_X1 U416 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U417 ( .A1(n608), .A2(n434), .ZN(n629) );
  INV_X1 U418 ( .A(KEYINPUT44), .ZN(n434) );
  XNOR2_X1 U419 ( .A(n398), .B(KEYINPUT81), .ZN(n452) );
  OR2_X1 U420 ( .A1(n593), .A2(n399), .ZN(n398) );
  NAND2_X1 U421 ( .A1(G953), .A2(n442), .ZN(n441) );
  XNOR2_X1 U422 ( .A(n489), .B(n490), .ZN(n380) );
  XNOR2_X1 U423 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n489) );
  XNOR2_X1 U424 ( .A(n735), .B(n458), .ZN(n525) );
  XNOR2_X1 U425 ( .A(n511), .B(n459), .ZN(n458) );
  INV_X1 U426 ( .A(KEYINPUT74), .ZN(n459) );
  NAND2_X1 U427 ( .A1(n375), .A2(n374), .ZN(n436) );
  AND2_X1 U428 ( .A1(n753), .A2(n589), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n376), .B(n582), .ZN(n375) );
  AND2_X1 U430 ( .A1(n577), .A2(n665), .ZN(n372) );
  NOR2_X1 U431 ( .A1(n612), .A2(KEYINPUT28), .ZN(n395) );
  INV_X1 U432 ( .A(n576), .ZN(n396) );
  NAND2_X1 U433 ( .A1(n612), .A2(KEYINPUT28), .ZN(n391) );
  XNOR2_X1 U434 ( .A(G902), .B(KEYINPUT15), .ZN(n635) );
  XNOR2_X1 U435 ( .A(n501), .B(KEYINPUT21), .ZN(n691) );
  XNOR2_X1 U436 ( .A(G107), .B(G122), .ZN(n516) );
  NOR2_X1 U437 ( .A1(n561), .A2(n568), .ZN(n562) );
  INV_X1 U438 ( .A(KEYINPUT34), .ZN(n384) );
  NAND2_X1 U439 ( .A1(n383), .A2(n435), .ZN(n688) );
  INV_X1 U440 ( .A(n691), .ZN(n435) );
  INV_X1 U441 ( .A(KEYINPUT1), .ZN(n579) );
  XNOR2_X1 U442 ( .A(n371), .B(n507), .ZN(n505) );
  XNOR2_X1 U443 ( .A(n382), .B(n743), .ZN(n642) );
  XNOR2_X1 U444 ( .A(n482), .B(n481), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n492), .B(KEYINPUT97), .ZN(n481) );
  XNOR2_X1 U446 ( .A(n496), .B(n495), .ZN(n482) );
  NAND2_X1 U447 ( .A1(n414), .A2(n366), .ZN(n638) );
  NAND2_X1 U448 ( .A1(n658), .A2(KEYINPUT47), .ZN(n463) );
  AND2_X1 U449 ( .A1(n450), .A2(n449), .ZN(n448) );
  NAND2_X1 U450 ( .A1(n691), .A2(n451), .ZN(n449) );
  INV_X1 U451 ( .A(G900), .ZN(n442) );
  INV_X1 U452 ( .A(KEYINPUT48), .ZN(n582) );
  INV_X1 U453 ( .A(KEYINPUT86), .ZN(n454) );
  XNOR2_X1 U454 ( .A(n443), .B(KEYINPUT92), .ZN(n591) );
  XNOR2_X1 U455 ( .A(n539), .B(n429), .ZN(n541) );
  XNOR2_X1 U456 ( .A(n540), .B(n430), .ZN(n429) );
  INV_X1 U457 ( .A(KEYINPUT103), .ZN(n430) );
  XNOR2_X1 U458 ( .A(G140), .B(G122), .ZN(n535) );
  XOR2_X1 U459 ( .A(G143), .B(G104), .Z(n536) );
  NOR2_X1 U460 ( .A1(G953), .A2(G237), .ZN(n543) );
  XNOR2_X1 U461 ( .A(KEYINPUT4), .B(G131), .ZN(n488) );
  XNOR2_X1 U462 ( .A(n521), .B(KEYINPUT10), .ZN(n544) );
  XOR2_X1 U463 ( .A(G137), .B(G140), .Z(n506) );
  XNOR2_X1 U464 ( .A(n388), .B(n353), .ZN(n387) );
  NAND2_X1 U465 ( .A1(n425), .A2(G227), .ZN(n388) );
  XOR2_X1 U466 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n518) );
  INV_X1 U467 ( .A(KEYINPUT4), .ZN(n517) );
  XNOR2_X1 U468 ( .A(n389), .B(KEYINPUT14), .ZN(n503) );
  NAND2_X1 U469 ( .A1(G234), .A2(G237), .ZN(n389) );
  OR2_X1 U470 ( .A1(G237), .A2(G902), .ZN(n526) );
  XNOR2_X1 U471 ( .A(n483), .B(n469), .ZN(n468) );
  XNOR2_X1 U472 ( .A(G116), .B(KEYINPUT99), .ZN(n483) );
  XNOR2_X1 U473 ( .A(KEYINPUT100), .B(KEYINPUT5), .ZN(n469) );
  BUF_X1 U474 ( .A(n672), .Z(n744) );
  XNOR2_X1 U475 ( .A(n373), .B(G119), .ZN(n515) );
  XNOR2_X1 U476 ( .A(G113), .B(KEYINPUT3), .ZN(n373) );
  XNOR2_X1 U477 ( .A(G104), .B(KEYINPUT78), .ZN(n508) );
  BUF_X1 U478 ( .A(n673), .Z(n732) );
  XNOR2_X1 U479 ( .A(G110), .B(KEYINPUT94), .ZN(n493) );
  XNOR2_X1 U480 ( .A(n672), .B(KEYINPUT79), .ZN(n460) );
  XNOR2_X1 U481 ( .A(n507), .B(n457), .ZN(n721) );
  XNOR2_X1 U482 ( .A(n525), .B(n385), .ZN(n457) );
  XNOR2_X1 U483 ( .A(n387), .B(n386), .ZN(n385) );
  INV_X1 U484 ( .A(n506), .ZN(n386) );
  AND2_X1 U485 ( .A1(n673), .A2(n472), .ZN(n677) );
  INV_X1 U486 ( .A(KEYINPUT2), .ZN(n473) );
  INV_X1 U487 ( .A(KEYINPUT19), .ZN(n470) );
  NAND2_X1 U488 ( .A1(n391), .A2(n610), .ZN(n390) );
  NAND2_X1 U489 ( .A1(n352), .A2(n362), .ZN(n561) );
  XNOR2_X1 U490 ( .A(n599), .B(KEYINPUT75), .ZN(n476) );
  XNOR2_X1 U491 ( .A(G475), .B(n550), .ZN(n566) );
  XNOR2_X1 U492 ( .A(n432), .B(n531), .ZN(n737) );
  XNOR2_X1 U493 ( .A(n515), .B(KEYINPUT16), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n532), .B(n419), .ZN(n727) );
  XNOR2_X1 U495 ( .A(n533), .B(n355), .ZN(n419) );
  NAND2_X1 U496 ( .A1(n725), .A2(G475), .ZN(n480) );
  XNOR2_X1 U497 ( .A(n587), .B(KEYINPUT107), .ZN(n753) );
  INV_X1 U498 ( .A(n402), .ZN(n587) );
  XNOR2_X1 U499 ( .A(n581), .B(KEYINPUT111), .ZN(n754) );
  INV_X1 U500 ( .A(KEYINPUT35), .ZN(n456) );
  NAND2_X1 U501 ( .A1(n623), .A2(n600), .ZN(n601) );
  NOR2_X1 U502 ( .A1(n383), .A2(n689), .ZN(n600) );
  NOR2_X1 U503 ( .A1(n615), .A2(n614), .ZN(n653) );
  NAND2_X1 U504 ( .A1(n424), .A2(n423), .ZN(n406) );
  XNOR2_X1 U505 ( .A(n640), .B(n365), .ZN(n424) );
  NAND2_X1 U506 ( .A1(n412), .A2(n423), .ZN(n407) );
  XNOR2_X1 U507 ( .A(n641), .B(n413), .ZN(n412) );
  INV_X1 U508 ( .A(n642), .ZN(n413) );
  INV_X1 U509 ( .A(KEYINPUT122), .ZN(n408) );
  INV_X1 U510 ( .A(KEYINPUT56), .ZN(n410) );
  XOR2_X1 U511 ( .A(G107), .B(KEYINPUT80), .Z(n353) );
  NAND2_X1 U512 ( .A1(n555), .A2(n403), .ZN(n354) );
  XNOR2_X1 U513 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n355) );
  AND2_X1 U514 ( .A1(n418), .A2(n417), .ZN(n356) );
  XOR2_X1 U515 ( .A(G128), .B(G119), .Z(n357) );
  AND2_X1 U516 ( .A1(n610), .A2(n552), .ZN(n358) );
  NOR2_X1 U517 ( .A1(KEYINPUT71), .A2(n683), .ZN(n359) );
  INV_X1 U518 ( .A(n404), .ZN(n623) );
  NAND2_X1 U519 ( .A1(n405), .A2(n605), .ZN(n404) );
  XOR2_X1 U520 ( .A(n499), .B(KEYINPUT25), .Z(n360) );
  AND2_X1 U521 ( .A1(G210), .A2(n526), .ZN(n361) );
  AND2_X1 U522 ( .A1(n358), .A2(n383), .ZN(n362) );
  XOR2_X1 U523 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n363) );
  XOR2_X1 U524 ( .A(n645), .B(n644), .Z(n364) );
  XOR2_X1 U525 ( .A(n505), .B(KEYINPUT62), .Z(n365) );
  XNOR2_X1 U526 ( .A(KEYINPUT66), .B(n637), .ZN(n366) );
  XOR2_X1 U527 ( .A(n723), .B(n722), .Z(n367) );
  XOR2_X1 U528 ( .A(n719), .B(n718), .Z(n368) );
  NOR2_X1 U529 ( .A1(G952), .A2(n425), .ZN(n729) );
  INV_X1 U530 ( .A(n729), .ZN(n423) );
  XOR2_X1 U531 ( .A(n646), .B(KEYINPUT67), .Z(n369) );
  XNOR2_X2 U532 ( .A(n578), .B(n470), .ZN(n431) );
  NAND2_X1 U533 ( .A1(n403), .A2(n678), .ZN(n578) );
  XNOR2_X2 U534 ( .A(n370), .B(G472), .ZN(n695) );
  XNOR2_X1 U535 ( .A(n486), .B(n487), .ZN(n371) );
  NAND2_X1 U536 ( .A1(n372), .A2(n678), .ZN(n583) );
  XNOR2_X1 U537 ( .A(n372), .B(KEYINPUT110), .ZN(n418) );
  XNOR2_X2 U538 ( .A(n436), .B(n634), .ZN(n672) );
  XNOR2_X2 U539 ( .A(n377), .B(n456), .ZN(n608) );
  NAND2_X1 U540 ( .A1(n378), .A2(n607), .ZN(n377) );
  XNOR2_X1 U541 ( .A(n379), .B(n384), .ZN(n378) );
  NAND2_X1 U542 ( .A1(n380), .A2(G221), .ZN(n496) );
  NAND2_X1 U543 ( .A1(n380), .A2(G217), .ZN(n533) );
  NOR2_X1 U544 ( .A1(n475), .A2(n383), .ZN(n474) );
  NAND2_X1 U545 ( .A1(n503), .A2(G902), .ZN(n443) );
  NAND2_X1 U546 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U547 ( .A1(n576), .A2(KEYINPUT28), .ZN(n393) );
  NAND2_X1 U548 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X2 U549 ( .A(n504), .B(n397), .ZN(n576) );
  INV_X1 U550 ( .A(KEYINPUT72), .ZN(n397) );
  NOR2_X1 U551 ( .A1(n591), .A2(n441), .ZN(n399) );
  AND2_X2 U552 ( .A1(n401), .A2(n400), .ZN(n630) );
  INV_X1 U553 ( .A(n656), .ZN(n400) );
  XNOR2_X1 U554 ( .A(n401), .B(G119), .ZN(G21) );
  XNOR2_X2 U555 ( .A(n601), .B(n363), .ZN(n401) );
  XNOR2_X1 U556 ( .A(n403), .B(KEYINPUT38), .ZN(n568) );
  OR2_X1 U557 ( .A1(n586), .A2(n403), .ZN(n402) );
  XNOR2_X2 U558 ( .A(n471), .B(n361), .ZN(n403) );
  NAND2_X1 U559 ( .A1(n405), .A2(n474), .ZN(n602) );
  XNOR2_X1 U560 ( .A(n406), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U561 ( .A(n407), .B(KEYINPUT125), .ZN(G66) );
  XNOR2_X1 U562 ( .A(n409), .B(n408), .ZN(G54) );
  NAND2_X1 U563 ( .A1(n422), .A2(n423), .ZN(n409) );
  XNOR2_X1 U564 ( .A(n411), .B(n410), .ZN(G51) );
  NAND2_X1 U565 ( .A1(n421), .A2(n423), .ZN(n411) );
  NAND2_X1 U566 ( .A1(n461), .A2(n460), .ZN(n414) );
  XNOR2_X2 U567 ( .A(n415), .B(G101), .ZN(n511) );
  NOR2_X2 U568 ( .A1(n570), .A2(n711), .ZN(n572) );
  XNOR2_X2 U569 ( .A(n514), .B(KEYINPUT108), .ZN(n570) );
  INV_X1 U570 ( .A(n578), .ZN(n417) );
  XNOR2_X1 U571 ( .A(n724), .B(n367), .ZN(n422) );
  XNOR2_X1 U572 ( .A(n720), .B(n368), .ZN(n421) );
  XNOR2_X1 U573 ( .A(n525), .B(n524), .ZN(n433) );
  XNOR2_X1 U574 ( .A(n433), .B(n737), .ZN(n717) );
  NAND2_X1 U575 ( .A1(n628), .A2(n627), .ZN(n455) );
  NAND2_X1 U576 ( .A1(n447), .A2(n446), .ZN(n445) );
  NAND2_X1 U577 ( .A1(n426), .A2(n462), .ZN(n438) );
  NOR2_X2 U578 ( .A1(n570), .A2(n431), .ZN(n662) );
  XNOR2_X1 U579 ( .A(n515), .B(n468), .ZN(n485) );
  NAND2_X1 U580 ( .A1(n695), .A2(n678), .ZN(n427) );
  NAND2_X1 U581 ( .A1(n759), .A2(n757), .ZN(n574) );
  NOR2_X2 U582 ( .A1(n431), .A2(n594), .ZN(n596) );
  INV_X1 U583 ( .A(n608), .ZN(n756) );
  INV_X1 U584 ( .A(n553), .ZN(n692) );
  OR2_X2 U585 ( .A1(n689), .A2(n688), .ZN(n617) );
  NOR2_X1 U586 ( .A1(n436), .A2(n473), .ZN(n472) );
  INV_X1 U587 ( .A(n754), .ZN(n440) );
  NOR2_X1 U588 ( .A1(n452), .A2(n691), .ZN(n552) );
  NOR2_X2 U589 ( .A1(n553), .A2(n444), .ZN(n504) );
  NOR2_X1 U590 ( .A1(n691), .A2(n451), .ZN(n446) );
  INV_X1 U591 ( .A(n452), .ZN(n447) );
  NAND2_X1 U592 ( .A1(n452), .A2(n451), .ZN(n450) );
  INV_X1 U593 ( .A(KEYINPUT73), .ZN(n451) );
  NAND2_X1 U594 ( .A1(n463), .A2(n556), .ZN(n462) );
  INV_X1 U595 ( .A(n662), .ZN(n658) );
  NAND2_X1 U596 ( .A1(n662), .A2(n465), .ZN(n464) );
  NAND2_X1 U597 ( .A1(n467), .A2(n560), .ZN(n466) );
  NAND2_X1 U598 ( .A1(n662), .A2(n359), .ZN(n467) );
  NAND2_X1 U599 ( .A1(n717), .A2(n635), .ZN(n471) );
  INV_X1 U600 ( .A(n612), .ZN(n475) );
  INV_X1 U601 ( .A(n635), .ZN(n477) );
  XNOR2_X1 U602 ( .A(n478), .B(n369), .ZN(G60) );
  XNOR2_X1 U603 ( .A(n574), .B(n573), .ZN(n575) );
  INV_X1 U604 ( .A(n647), .ZN(n625) );
  XNOR2_X1 U605 ( .A(n519), .B(n518), .ZN(n523) );
  INV_X1 U606 ( .A(n670), .ZN(n589) );
  INV_X1 U607 ( .A(G469), .ZN(n512) );
  XNOR2_X1 U608 ( .A(n511), .B(G137), .ZN(n487) );
  NAND2_X1 U609 ( .A1(n543), .A2(G210), .ZN(n484) );
  XNOR2_X1 U610 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X2 U611 ( .A(G128), .B(G143), .Z(n520) );
  NAND2_X1 U612 ( .A1(n745), .A2(G234), .ZN(n490) );
  XNOR2_X1 U613 ( .A(KEYINPUT96), .B(KEYINPUT24), .ZN(n491) );
  XNOR2_X1 U614 ( .A(n357), .B(n491), .ZN(n492) );
  XOR2_X1 U615 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n494) );
  XNOR2_X1 U616 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U617 ( .A(n506), .B(n544), .ZN(n743) );
  NAND2_X1 U618 ( .A1(n635), .A2(G234), .ZN(n498) );
  XNOR2_X1 U619 ( .A(n498), .B(n497), .ZN(n500) );
  NAND2_X1 U620 ( .A1(G217), .A2(n500), .ZN(n499) );
  NAND2_X1 U621 ( .A1(n500), .A2(G221), .ZN(n501) );
  NAND2_X1 U622 ( .A1(G952), .A2(n503), .ZN(n707) );
  XNOR2_X1 U623 ( .A(n502), .B(KEYINPUT90), .ZN(n593) );
  INV_X1 U624 ( .A(n508), .ZN(n510) );
  XNOR2_X1 U625 ( .A(G110), .B(KEYINPUT89), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n510), .B(n509), .ZN(n735) );
  NOR2_X1 U627 ( .A1(G902), .A2(n721), .ZN(n513) );
  XNOR2_X1 U628 ( .A(n516), .B(G116), .ZN(n531) );
  XNOR2_X1 U629 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U630 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U631 ( .A1(G214), .A2(n526), .ZN(n678) );
  INV_X1 U632 ( .A(KEYINPUT71), .ZN(n527) );
  INV_X1 U633 ( .A(KEYINPUT47), .ZN(n551) );
  AND2_X1 U634 ( .A1(n527), .A2(n551), .ZN(n528) );
  INV_X1 U635 ( .A(n529), .ZN(n530) );
  XNOR2_X1 U636 ( .A(n531), .B(n530), .ZN(n532) );
  NOR2_X1 U637 ( .A1(G902), .A2(n727), .ZN(n534) );
  XOR2_X1 U638 ( .A(G478), .B(n534), .Z(n565) );
  XNOR2_X1 U639 ( .A(n536), .B(n535), .ZN(n542) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(KEYINPUT104), .Z(n538) );
  XNOR2_X1 U641 ( .A(KEYINPUT12), .B(KEYINPUT102), .ZN(n537) );
  XNOR2_X1 U642 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U643 ( .A(n542), .B(n541), .ZN(n547) );
  NAND2_X1 U644 ( .A1(n543), .A2(G214), .ZN(n545) );
  XNOR2_X1 U645 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n547), .B(n546), .ZN(n643) );
  NOR2_X1 U647 ( .A1(G902), .A2(n643), .ZN(n549) );
  XNOR2_X1 U648 ( .A(KEYINPUT105), .B(KEYINPUT13), .ZN(n548) );
  XNOR2_X1 U649 ( .A(n549), .B(n548), .ZN(n550) );
  INV_X1 U650 ( .A(n665), .ZN(n563) );
  NAND2_X1 U651 ( .A1(n565), .A2(n566), .ZN(n659) );
  NAND2_X1 U652 ( .A1(n563), .A2(n659), .ZN(n559) );
  INV_X1 U653 ( .A(n566), .ZN(n554) );
  NAND2_X1 U654 ( .A1(n565), .A2(n554), .ZN(n604) );
  NOR2_X1 U655 ( .A1(n561), .A2(n604), .ZN(n555) );
  NAND2_X1 U656 ( .A1(n354), .A2(KEYINPUT82), .ZN(n556) );
  INV_X1 U657 ( .A(KEYINPUT82), .ZN(n557) );
  NAND2_X1 U658 ( .A1(n559), .A2(n557), .ZN(n558) );
  AND2_X1 U659 ( .A1(n558), .A2(KEYINPUT47), .ZN(n560) );
  INV_X1 U660 ( .A(n559), .ZN(n683) );
  XNOR2_X1 U661 ( .A(n562), .B(KEYINPUT39), .ZN(n588) );
  INV_X1 U662 ( .A(n565), .ZN(n567) );
  NAND2_X1 U663 ( .A1(n567), .A2(n566), .ZN(n681) );
  INV_X1 U664 ( .A(n568), .ZN(n679) );
  NAND2_X1 U665 ( .A1(n679), .A2(n678), .ZN(n682) );
  NOR2_X1 U666 ( .A1(n681), .A2(n682), .ZN(n569) );
  XNOR2_X1 U667 ( .A(n569), .B(KEYINPUT41), .ZN(n711) );
  XNOR2_X1 U668 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n571) );
  XNOR2_X1 U669 ( .A(n572), .B(n571), .ZN(n757) );
  XOR2_X1 U670 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n573) );
  XNOR2_X1 U671 ( .A(n695), .B(KEYINPUT6), .ZN(n605) );
  NOR2_X1 U672 ( .A1(n576), .A2(n605), .ZN(n577) );
  XNOR2_X1 U673 ( .A(KEYINPUT36), .B(n356), .ZN(n580) );
  INV_X1 U674 ( .A(n689), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n580), .A2(n603), .ZN(n581) );
  XNOR2_X1 U676 ( .A(KEYINPUT106), .B(n583), .ZN(n584) );
  NOR2_X1 U677 ( .A1(n603), .A2(n584), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n585), .B(KEYINPUT43), .ZN(n586) );
  NOR2_X1 U679 ( .A1(n588), .A2(n659), .ZN(n670) );
  NOR2_X1 U680 ( .A1(G898), .A2(n425), .ZN(n590) );
  XNOR2_X1 U681 ( .A(KEYINPUT91), .B(n590), .ZN(n739) );
  NOR2_X1 U682 ( .A1(n591), .A2(n739), .ZN(n592) );
  NOR2_X1 U683 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X2 U684 ( .A(n596), .B(n595), .ZN(n616) );
  NOR2_X1 U685 ( .A1(n681), .A2(n691), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n616), .A2(n597), .ZN(n598) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n599) );
  NOR2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n656) );
  INV_X1 U689 ( .A(n604), .ZN(n607) );
  NOR2_X1 U690 ( .A1(n617), .A2(n605), .ZN(n606) );
  XNOR2_X1 U691 ( .A(KEYINPUT33), .B(n606), .ZN(n710) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT93), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n630), .A2(n608), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n609), .A2(KEYINPUT44), .ZN(n628) );
  INV_X1 U695 ( .A(n610), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n611), .A2(n688), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U698 ( .A(n616), .ZN(n619) );
  INV_X1 U699 ( .A(n617), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n695), .A2(n618), .ZN(n698) );
  NOR2_X1 U701 ( .A1(n619), .A2(n698), .ZN(n621) );
  XNOR2_X1 U702 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n621), .B(n620), .ZN(n668) );
  NOR2_X1 U704 ( .A1(n653), .A2(n668), .ZN(n622) );
  NOR2_X1 U705 ( .A1(n683), .A2(n622), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n692), .A2(n404), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n689), .A2(n624), .ZN(n647) );
  XNOR2_X1 U708 ( .A(KEYINPUT70), .B(n629), .ZN(n632) );
  XOR2_X1 U709 ( .A(n630), .B(KEYINPUT87), .Z(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  INV_X1 U711 ( .A(n677), .ZN(n639) );
  XOR2_X1 U712 ( .A(n635), .B(KEYINPUT84), .Z(n636) );
  NAND2_X1 U713 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G472), .A2(n725), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G217), .A2(n725), .ZN(n641) );
  XNOR2_X1 U716 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT123), .ZN(n644) );
  INV_X1 U718 ( .A(KEYINPUT60), .ZN(n646) );
  XNOR2_X1 U719 ( .A(G101), .B(n647), .ZN(G3) );
  NAND2_X1 U720 ( .A1(n653), .A2(n665), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(KEYINPUT112), .ZN(n649) );
  XNOR2_X1 U722 ( .A(G104), .B(n649), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n651) );
  XNOR2_X1 U724 ( .A(G107), .B(KEYINPUT113), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U726 ( .A(KEYINPUT26), .B(n652), .Z(n655) );
  INV_X1 U727 ( .A(n659), .ZN(n667) );
  NAND2_X1 U728 ( .A1(n653), .A2(n667), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(G9) );
  XNOR2_X1 U730 ( .A(G110), .B(n656), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(KEYINPUT115), .ZN(G12) );
  NOR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U733 ( .A(G128), .B(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(G30) );
  XNOR2_X1 U735 ( .A(G143), .B(n354), .ZN(G45) );
  NAND2_X1 U736 ( .A1(n662), .A2(n665), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(KEYINPUT116), .ZN(n664) );
  XNOR2_X1 U738 ( .A(G146), .B(n664), .ZN(G48) );
  NAND2_X1 U739 ( .A1(n668), .A2(n665), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n666), .B(G113), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(G116), .ZN(G18) );
  XNOR2_X1 U743 ( .A(G134), .B(n670), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT117), .ZN(G36) );
  INV_X1 U745 ( .A(n732), .ZN(n674) );
  NOR2_X1 U746 ( .A1(n744), .A2(n674), .ZN(n675) );
  NOR2_X1 U747 ( .A1(KEYINPUT2), .A2(n675), .ZN(n676) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n709) );
  NOR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n686), .A2(n710), .ZN(n687) );
  XOR2_X1 U754 ( .A(KEYINPUT119), .B(n687), .Z(n704) );
  NAND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT50), .ZN(n697) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U758 ( .A(KEYINPUT49), .B(n693), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n475), .A2(n694), .ZN(n696) );
  NAND2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U762 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n711), .A2(n701), .ZN(n702) );
  XNOR2_X1 U764 ( .A(KEYINPUT118), .B(n702), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U766 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U770 ( .A(KEYINPUT120), .B(n712), .Z(n713) );
  NAND2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n715), .A2(G953), .ZN(n716) );
  XNOR2_X1 U773 ( .A(n716), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U774 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n717), .B(KEYINPUT88), .ZN(n718) );
  NAND2_X1 U776 ( .A1(n725), .A2(G210), .ZN(n720) );
  XNOR2_X1 U777 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n723) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT57), .ZN(n722) );
  NAND2_X1 U779 ( .A1(n725), .A2(G469), .ZN(n724) );
  NAND2_X1 U780 ( .A1(G478), .A2(n725), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n729), .A2(n728), .ZN(G63) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n731), .A2(G898), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n732), .A2(n425), .ZN(n733) );
  NAND2_X1 U787 ( .A1(n734), .A2(n733), .ZN(n741) );
  XOR2_X1 U788 ( .A(n735), .B(G101), .Z(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U791 ( .A(n741), .B(n740), .Z(G69) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(n748) );
  XNOR2_X1 U793 ( .A(n748), .B(n744), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(n425), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n747), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U796 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G953), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n752), .A2(n751), .ZN(G72) );
  XNOR2_X1 U800 ( .A(G140), .B(n753), .ZN(G42) );
  XNOR2_X1 U801 ( .A(n754), .B(G125), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n755), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U803 ( .A(n756), .B(G122), .Z(G24) );
  XOR2_X1 U804 ( .A(G137), .B(n757), .Z(n758) );
  XNOR2_X1 U805 ( .A(KEYINPUT127), .B(n758), .ZN(G39) );
  XNOR2_X1 U806 ( .A(G131), .B(n759), .ZN(G33) );
endmodule

