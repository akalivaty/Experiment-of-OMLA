//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n203), .A2(G1gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n206), .A2(new_n207), .A3(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  XOR2_X1   g008(.A(G15gat), .B(G22gat), .Z(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n203), .A2(new_n205), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n202), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(G8gat), .B1(new_n206), .B2(new_n207), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n209), .A3(new_n212), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT90), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT15), .B1(new_n218), .B2(KEYINPUT89), .ZN(new_n219));
  OR2_X1    g018(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G50gat), .ZN(new_n227));
  INV_X1    g026(.A(G50gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G43gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G29gat), .ZN(new_n231));
  INV_X1    g030(.A(G36gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT14), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT14), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G29gat), .B2(G36gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n219), .A2(new_n223), .A3(new_n230), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n232), .B1(new_n220), .B2(new_n221), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n235), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT15), .B(new_n218), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n237), .B2(new_n241), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n214), .B(new_n217), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n208), .A2(new_n213), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n237), .A2(new_n241), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n249), .A4(new_n245), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(new_n241), .A3(new_n237), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n245), .B(KEYINPUT13), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G169gat), .B(G197gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT12), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n252), .A2(new_n253), .A3(new_n257), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT91), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n250), .A2(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT91), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n253), .A4(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n253), .ZN(new_n270));
  INV_X1    g069(.A(new_n263), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G22gat), .ZN(new_n275));
  XOR2_X1   g074(.A(G141gat), .B(G148gat), .Z(new_n276));
  INV_X1    g075(.A(G155gat), .ZN(new_n277));
  INV_X1    g076(.A(G162gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT2), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G155gat), .B(G162gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT29), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT73), .ZN(new_n286));
  XOR2_X1   g085(.A(G197gat), .B(G204gat), .Z(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT72), .B(G211gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G218gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n286), .B(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G228gat), .A2(G233gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT3), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n282), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n293), .A2(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(KEYINPUT77), .ZN(new_n300));
  INV_X1    g099(.A(new_n292), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n291), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(KEYINPUT76), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(KEYINPUT29), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT3), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n299), .B(new_n300), .C1(new_n306), .C2(new_n282), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n294), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n307), .B2(new_n294), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n275), .B(new_n298), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT79), .ZN(new_n313));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT31), .B(G50gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n298), .B1(new_n310), .B2(new_n311), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G22gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n312), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n322));
  NOR2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT64), .B(G190gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(KEYINPUT28), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n332), .A2(new_n329), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n334), .A2(KEYINPUT28), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n328), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT24), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT24), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(G183gat), .B2(G190gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n325), .B1(new_n323), .B2(KEYINPUT23), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(KEYINPUT23), .B2(new_n323), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n337), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT65), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n341), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(KEYINPUT65), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT25), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n355));
  XNOR2_X1  g154(.A(G127gat), .B(G134gat), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(G120gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT1), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT68), .B(G113gat), .Z(new_n360));
  OAI211_X1 g159(.A(new_n356), .B(new_n359), .C1(new_n360), .C2(new_n358), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n356), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n365));
  NAND2_X1  g164(.A1(G113gat), .A2(G120gat), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n364), .A2(new_n365), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n365), .B2(new_n364), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n355), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n353), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n363), .A2(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT70), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n322), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G71gat), .B(G99gat), .Z(new_n380));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n375), .A2(new_n377), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n379), .B(new_n382), .C1(KEYINPUT33), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(KEYINPUT33), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n378), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n378), .B2(new_n386), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n370), .A2(new_n376), .A3(new_n374), .A4(new_n373), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT34), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n384), .B(new_n392), .C1(new_n388), .C2(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n319), .A2(new_n396), .A3(new_n312), .A4(new_n316), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n321), .A2(new_n394), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n354), .B2(KEYINPUT29), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n371), .A2(G226gat), .A3(G233gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n301), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n292), .A3(new_n404), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n401), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n407), .A3(new_n401), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(KEYINPUT30), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n407), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n401), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n369), .A2(new_n282), .ZN(new_n418));
  INV_X1    g217(.A(new_n282), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n372), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n282), .B(new_n283), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n425), .A2(new_n369), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n372), .A2(new_n419), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .A4(new_n422), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n418), .B(KEYINPUT4), .C1(new_n369), .C2(new_n425), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n424), .A2(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G57gat), .B(G85gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT6), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT6), .B1(new_n436), .B2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n445), .B2(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n416), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT35), .B1(new_n398), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n397), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n313), .A2(new_n316), .B1(new_n319), .B2(new_n312), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n395), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n378), .A2(new_n386), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n387), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n392), .B1(new_n455), .B2(new_n384), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n416), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n441), .B(KEYINPUT80), .Z(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n436), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n431), .A2(new_n424), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n434), .A2(new_n435), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n461), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(KEYINPUT83), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n444), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n443), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n451), .A2(new_n457), .A3(new_n459), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n448), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT38), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n401), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n408), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n407), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n403), .A2(KEYINPUT85), .A3(new_n292), .A4(new_n404), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n406), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n480), .A2(KEYINPUT86), .A3(KEYINPUT37), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT86), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n473), .B(new_n476), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n413), .A2(new_n474), .B1(new_n408), .B2(new_n475), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n484), .A2(KEYINPUT38), .B1(new_n413), .B2(new_n401), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n483), .A2(new_n485), .A3(new_n443), .A4(new_n469), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n411), .A2(new_n415), .A3(new_n468), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n418), .A2(new_n422), .A3(new_n420), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT39), .B(new_n488), .C1(new_n434), .C2(new_n422), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT81), .B(KEYINPUT39), .Z(new_n490));
  NAND4_X1  g289(.A1(new_n432), .A2(new_n423), .A3(new_n433), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n461), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT82), .B1(new_n491), .B2(new_n461), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT40), .B(new_n489), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT40), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n493), .A2(new_n494), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n432), .A2(new_n423), .A3(new_n433), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n500), .A2(KEYINPUT39), .A3(new_n488), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n503), .A3(new_n451), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n452), .B2(new_n456), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n394), .A2(KEYINPUT36), .A3(new_n395), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n321), .A2(new_n397), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n447), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n274), .B1(new_n472), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT93), .B1(new_n513), .B2(KEYINPUT9), .ZN(new_n514));
  INV_X1    g313(.A(G57gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G64gat), .ZN(new_n516));
  INV_X1    g315(.A(G64gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G57gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n516), .A2(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n526), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n514), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G127gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n247), .B1(KEYINPUT21), .B2(new_n534), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G155gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G183gat), .B(G211gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n541), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n548), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n547), .ZN(new_n557));
  NOR2_X1   g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n557), .A2(new_n558), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n560), .A2(KEYINPUT94), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT94), .B1(new_n560), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n248), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n242), .A2(new_n243), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n570), .B(new_n572), .C1(new_n573), .C2(new_n569), .ZN(new_n574));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT95), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n574), .A2(new_n577), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n582), .A2(KEYINPUT96), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT97), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n584), .B2(new_n585), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n546), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n556), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n564), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n556), .A2(new_n559), .A3(new_n594), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n531), .A2(new_n514), .A3(new_n532), .ZN(new_n598));
  NAND2_X1  g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n524), .B1(new_n601), .B2(new_n526), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n531), .B2(new_n514), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n556), .A2(new_n559), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n530), .B(new_n533), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT10), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n530), .B2(new_n533), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n605), .B2(new_n606), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n560), .A2(KEYINPUT94), .A3(new_n566), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n593), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n593), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n604), .A2(new_n607), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT99), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n616), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n616), .B2(new_n618), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n592), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n512), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n446), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT100), .B(G1gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1324gat));
  INV_X1    g431(.A(new_n628), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT16), .B(G8gat), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n633), .A2(new_n416), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n209), .B1(new_n628), .B2(new_n458), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT42), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(KEYINPUT42), .B2(new_n635), .ZN(G1325gat));
  NOR3_X1   g437(.A1(new_n452), .A2(new_n456), .A3(new_n505), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT36), .B1(new_n394), .B2(new_n395), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT101), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n506), .A2(new_n642), .A3(new_n507), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G15gat), .B1(new_n633), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n457), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n633), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n628), .A2(new_n509), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT102), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n546), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n625), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n591), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n512), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n656), .A2(new_n629), .A3(new_n220), .A4(new_n221), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n641), .A2(new_n510), .A3(new_n504), .A4(new_n643), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n472), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n590), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n472), .A2(new_n511), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n591), .A2(new_n663), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n662), .A2(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n654), .A2(new_n274), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n222), .B1(new_n668), .B2(new_n446), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n659), .A2(new_n669), .ZN(G1328gat));
  NAND3_X1  g469(.A1(new_n656), .A2(new_n232), .A3(new_n458), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G36gat), .B1(new_n668), .B2(new_n416), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(KEYINPUT104), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  OAI21_X1  g478(.A(G43gat), .B1(new_n668), .B2(new_n644), .ZN(new_n680));
  NOR2_X1   g479(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n646), .A2(G43gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n656), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1330gat));
  NAND4_X1  g485(.A1(new_n666), .A2(G50gat), .A3(new_n509), .A4(new_n667), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT48), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n656), .A2(new_n509), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n228), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n687), .A2(new_n690), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(KEYINPUT48), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT107), .B(new_n688), .C1(new_n687), .C2(new_n690), .ZN(new_n697));
  OAI22_X1  g496(.A1(new_n692), .A2(new_n693), .B1(new_n696), .B2(new_n697), .ZN(G1331gat));
  NOR3_X1   g497(.A1(new_n592), .A2(new_n273), .A3(new_n625), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n661), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n629), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g501(.A1(new_n700), .A2(new_n458), .ZN(new_n703));
  NOR2_X1   g502(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n704));
  AND2_X1   g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n703), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT108), .ZN(G1333gat));
  INV_X1    g507(.A(new_n644), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n646), .A2(G71gat), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n710), .A2(G71gat), .B1(new_n700), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g512(.A1(new_n700), .A2(new_n509), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g514(.A1(new_n446), .A2(G85gat), .A3(new_n625), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n546), .A2(new_n273), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n661), .A2(KEYINPUT51), .A3(new_n590), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT110), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n661), .A2(new_n590), .A3(new_n717), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n591), .B1(new_n660), .B2(new_n472), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT51), .A4(new_n717), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(KEYINPUT111), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(KEYINPUT111), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n716), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n664), .A2(new_n665), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n717), .A2(new_n626), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT109), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n732), .C1(new_n723), .C2(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n446), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(G1336gat));
  OAI21_X1  g534(.A(G92gat), .B1(new_n733), .B2(new_n416), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n416), .A2(G92gat), .A3(new_n625), .ZN(new_n737));
  INV_X1    g536(.A(new_n718), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n723), .B2(new_n717), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT52), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n666), .A2(new_n743), .A3(new_n458), .A4(new_n732), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT112), .B1(new_n733), .B2(new_n416), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n745), .A3(G92gat), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT52), .B1(new_n726), .B2(new_n737), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n749), .B2(new_n750), .ZN(G1337gat));
  NOR3_X1   g550(.A1(new_n646), .A2(G99gat), .A3(new_n625), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT114), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n727), .B2(new_n728), .ZN(new_n754));
  OAI21_X1  g553(.A(G99gat), .B1(new_n733), .B2(new_n644), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1338gat));
  NOR3_X1   g555(.A1(new_n451), .A2(G106gat), .A3(new_n625), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n726), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  OAI21_X1  g558(.A(G106gat), .B1(new_n733), .B2(new_n451), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n762), .B(G106gat), .C1(new_n733), .C2(new_n451), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(KEYINPUT115), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n757), .B1(new_n738), .B2(new_n739), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n767), .B(new_n757), .C1(new_n738), .C2(new_n739), .ZN(new_n768));
  AND4_X1   g567(.A1(new_n763), .A2(new_n764), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n761), .B1(new_n769), .B2(new_n759), .ZN(G1339gat));
  NOR3_X1   g569(.A1(new_n592), .A2(new_n273), .A3(new_n626), .ZN(new_n771));
  INV_X1    g570(.A(new_n623), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n604), .A2(new_n607), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n609), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n617), .B1(new_n774), .B2(new_n614), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n614), .A2(new_n617), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT54), .B1(new_n776), .B2(new_n608), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n593), .B1(new_n569), .B2(new_n610), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT117), .B1(new_n782), .B2(new_n616), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT55), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n780), .B(new_n593), .C1(new_n608), .C2(new_n615), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786));
  INV_X1    g585(.A(new_n622), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n772), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n787), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT118), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n778), .B1(new_n775), .B2(new_n777), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n782), .A2(KEYINPUT117), .A3(new_n616), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT55), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n262), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n255), .A2(new_n256), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n244), .A2(new_n249), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(G229gat), .A3(G233gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n265), .B2(new_n268), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n800), .A2(new_n590), .A3(new_n806), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n805), .B(new_n625), .C1(new_n265), .C2(new_n268), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n800), .B2(new_n273), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(new_n590), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n546), .B1(new_n810), .B2(KEYINPUT119), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n807), .C1(new_n809), .C2(new_n590), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n771), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n446), .ZN(new_n815));
  INV_X1    g614(.A(new_n398), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n458), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n360), .A3(new_n273), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n814), .A2(new_n509), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n458), .A2(new_n446), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n457), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n274), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1340gat));
  NOR3_X1   g623(.A1(new_n822), .A2(new_n358), .A3(new_n625), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n626), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n358), .ZN(G1341gat));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n538), .A3(new_n546), .ZN(new_n828));
  OAI21_X1  g627(.A(G127gat), .B1(new_n822), .B2(new_n653), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1342gat));
  OR4_X1    g629(.A1(G134gat), .A2(new_n817), .A3(new_n458), .A4(new_n591), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n822), .B2(new_n591), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(G1343gat));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT120), .B(new_n836), .C1(new_n814), .C2(new_n451), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n795), .A2(new_n798), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n796), .B2(new_n797), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n623), .B1(new_n842), .B2(new_n795), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n273), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n806), .A2(new_n626), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n590), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND4_X1   g645(.A1(new_n590), .A2(new_n841), .A3(new_n806), .A4(new_n843), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT119), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n813), .A3(new_n653), .ZN(new_n849));
  INV_X1    g648(.A(new_n771), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n451), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n838), .B1(new_n851), .B2(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n810), .A2(new_n653), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(KEYINPUT57), .A3(new_n509), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n641), .A2(new_n643), .A3(new_n821), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n274), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n641), .A2(new_n509), .A3(new_n643), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n815), .A3(new_n416), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(G141gat), .A3(new_n274), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n856), .A2(KEYINPUT121), .A3(new_n857), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT121), .B1(new_n856), .B2(new_n857), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n866), .A2(new_n867), .A3(new_n274), .ZN(new_n868));
  INV_X1    g667(.A(G141gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT122), .B1(new_n870), .B2(KEYINPUT58), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n858), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n856), .A2(KEYINPUT121), .A3(new_n857), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n273), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n862), .B1(new_n875), .B2(G141gat), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n864), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n865), .B1(new_n871), .B2(new_n878), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n509), .A2(KEYINPUT57), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n451), .B1(new_n850), .B2(new_n853), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n814), .A2(new_n880), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(new_n857), .A3(new_n626), .ZN(new_n883));
  INV_X1    g682(.A(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT59), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n866), .A2(new_n867), .A3(new_n625), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n884), .A2(KEYINPUT59), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n861), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n884), .A3(new_n626), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1345gat));
  AOI21_X1  g690(.A(G155gat), .B1(new_n889), .B2(new_n546), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n866), .A2(new_n867), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n546), .A2(G155gat), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT123), .Z(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT124), .ZN(G1346gat));
  NOR3_X1   g696(.A1(new_n458), .A2(G162gat), .A3(new_n591), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n860), .A2(new_n815), .A3(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n866), .A2(new_n867), .A3(new_n591), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n278), .ZN(G1347gat));
  NOR3_X1   g700(.A1(new_n646), .A2(new_n629), .A3(new_n416), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n820), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n274), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n816), .A2(new_n458), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT125), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n814), .A2(new_n629), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n273), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n905), .B1(new_n911), .B2(new_n904), .ZN(G1348gat));
  OAI21_X1  g711(.A(G176gat), .B1(new_n903), .B2(new_n625), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n625), .A2(G176gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n909), .B2(new_n914), .ZN(G1349gat));
  INV_X1    g714(.A(new_n903), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n337), .B1(new_n916), .B2(new_n546), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n546), .A2(new_n331), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n903), .B2(new_n591), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT61), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n910), .A2(new_n332), .A3(new_n590), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1351gat));
  AND2_X1   g724(.A1(new_n860), .A2(new_n458), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n908), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n273), .ZN(new_n929));
  AND4_X1   g728(.A1(new_n446), .A2(new_n882), .A3(new_n458), .A4(new_n644), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n273), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  OR2_X1    g731(.A1(new_n625), .A2(G204gat), .ZN(new_n933));
  OR3_X1    g732(.A1(new_n927), .A2(KEYINPUT62), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n626), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G204gat), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT62), .B1(new_n927), .B2(new_n933), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(G1353gat));
  OR3_X1    g737(.A1(new_n927), .A2(new_n288), .A3(new_n653), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n930), .A2(new_n546), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n928), .B2(new_n590), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n590), .A2(G218gat), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT127), .Z(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n930), .B2(new_n946), .ZN(G1355gat));
endmodule


