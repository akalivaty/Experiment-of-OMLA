//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  OR2_X1    g001(.A1(KEYINPUT66), .A2(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT66), .A2(G119), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G116), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n187), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n187), .B1(new_n190), .B2(new_n192), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT30), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G128), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n202), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(G128), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n200), .A2(new_n206), .A3(G143), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(KEYINPUT65), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n201), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT64), .A2(G131), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT64), .A2(G131), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G137), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(G137), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n222), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n233), .B(new_n234), .C1(new_n205), .C2(new_n207), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT0), .A4(G128), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n226), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n198), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT65), .B1(new_n213), .B2(new_n214), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n209), .B(new_n202), .C1(new_n199), .C2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n243), .A2(new_n244), .B1(new_n199), .B2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n241), .B(new_n198), .C1(new_n246), .C2(new_n230), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n197), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(G953), .ZN(new_n250));
  INV_X1    g064(.A(G237), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(G210), .A3(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n241), .B(new_n196), .C1(new_n246), .C2(new_n230), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n249), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT31), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n241), .B1(new_n246), .B2(new_n230), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n197), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n264), .B2(new_n258), .ZN(new_n265));
  INV_X1    g079(.A(new_n258), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n256), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(KEYINPUT30), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n247), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n270), .B2(new_n197), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n257), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n260), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G472), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT32), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n275), .A4(new_n276), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n275), .A4(new_n276), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n196), .B1(new_n232), .B2(new_n241), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT28), .B1(new_n284), .B2(new_n266), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n264), .A2(new_n258), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n258), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT72), .B1(new_n258), .B2(new_n290), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n256), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n287), .A2(new_n289), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n276), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n299), .A3(new_n276), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n271), .A2(new_n256), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n257), .B1(new_n265), .B2(new_n267), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G472), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n282), .A2(new_n283), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G125), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G140), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT16), .ZN(new_n312));
  OR3_X1    g126(.A1(new_n310), .A2(KEYINPUT16), .A3(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n206), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n313), .A3(G146), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G119), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n188), .A2(new_n189), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G128), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT24), .B(G110), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G110), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n324));
  AOI21_X1  g138(.A(G128), .B1(new_n188), .B2(new_n189), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n323), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n309), .A2(new_n311), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n206), .ZN(new_n331));
  AND4_X1   g145(.A1(new_n329), .A2(new_n309), .A3(new_n311), .A4(new_n206), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n316), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n323), .A3(new_n326), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n320), .A2(new_n321), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n250), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G137), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n328), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n322), .A2(new_n327), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n345), .A2(new_n346), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G217), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(G234), .B2(new_n276), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT74), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n341), .A2(new_n344), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n352), .A2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n307), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G214), .B1(G237), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G104), .ZN(new_n368));
  AOI21_X1  g182(.A(G107), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G104), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT81), .B(G101), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n371), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT77), .B(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(G107), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT81), .B1(new_n376), .B2(G101), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n370), .A3(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n383), .A2(new_n380), .A3(new_n370), .A4(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n366), .A2(new_n368), .A3(G107), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n379), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n190), .A2(KEYINPUT5), .A3(new_n192), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n188), .A2(new_n390), .A3(G116), .A4(new_n189), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n393));
  OAI211_X1 g207(.A(G113), .B(new_n389), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n378), .A2(new_n193), .A3(new_n388), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n387), .B1(new_n369), .B2(new_n380), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n383), .B1(new_n398), .B2(new_n370), .ZN(new_n399));
  INV_X1    g213(.A(new_n384), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n379), .A2(new_n385), .A3(KEYINPUT79), .A4(new_n387), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(G101), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n388), .A2(KEYINPUT4), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n197), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n395), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(new_n395), .C1(new_n406), .C2(new_n409), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT6), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n404), .A2(new_n405), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n197), .A3(new_n408), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n412), .B1(new_n418), .B2(new_n395), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n364), .B(new_n414), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n413), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n421), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n415), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n310), .B1(new_n235), .B2(new_n236), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n246), .B2(new_n310), .ZN(new_n425));
  INV_X1    g239(.A(G953), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G224), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n425), .B(new_n427), .Z(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G210), .B1(G237), .B2(G902), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT89), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n246), .A2(new_n310), .ZN(new_n434));
  INV_X1    g248(.A(new_n424), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(KEYINPUT7), .A3(new_n435), .A4(new_n427), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT87), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n425), .A2(new_n438), .A3(KEYINPUT7), .A4(new_n427), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n412), .B(KEYINPUT8), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n394), .A2(new_n193), .ZN(new_n442));
  OAI21_X1  g256(.A(G101), .B1(new_n369), .B2(new_n371), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n388), .A3(new_n372), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n378), .A2(new_n388), .B1(new_n394), .B2(new_n193), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n441), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n425), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n451));
  AOI22_X1  g265(.A1(KEYINPUT86), .A2(new_n451), .B1(new_n426), .B2(G224), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(KEYINPUT86), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n440), .A2(KEYINPUT88), .A3(new_n449), .A4(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n455), .A2(new_n415), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n446), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n395), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n458), .A2(new_n441), .B1(new_n450), .B2(new_n453), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT88), .B1(new_n459), .B2(new_n440), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n430), .A2(new_n433), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n428), .B1(new_n420), .B2(new_n422), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(new_n415), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n276), .B1(new_n465), .B2(new_n460), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n432), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n363), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n426), .A2(G952), .ZN(new_n469));
  INV_X1    g283(.A(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n251), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n276), .B(new_n250), .C1(G234), .C2(G237), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n426), .A2(KEYINPUT67), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G953), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n478), .A2(new_n480), .A3(G214), .A4(new_n251), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n204), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n250), .A2(G143), .A3(G214), .A4(new_n251), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n477), .B(new_n219), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT90), .B1(new_n484), .B2(new_n317), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(new_n219), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(KEYINPUT17), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n315), .A4(new_n316), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n483), .A3(new_n219), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n477), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n365), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n486), .A2(KEYINPUT18), .A3(G131), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT18), .A2(G131), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n483), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n331), .A2(new_n332), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n330), .A2(new_n206), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n497), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n494), .A2(new_n496), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT91), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n494), .A2(new_n505), .A3(new_n496), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n491), .A2(new_n492), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n330), .B(KEYINPUT19), .Z(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(new_n316), .C1(G146), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n496), .B1(new_n510), .B2(new_n502), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n511), .B1(new_n504), .B2(new_n506), .ZN(new_n517));
  INV_X1    g331(.A(new_n515), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT20), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n496), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n494), .A2(new_n502), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n504), .A2(new_n506), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G475), .B1(new_n523), .B2(G902), .ZN(new_n524));
  INV_X1    g338(.A(G478), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT9), .B(G234), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n527), .A2(new_n351), .A3(G953), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n191), .A2(G122), .ZN(new_n529));
  INV_X1    g343(.A(G122), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G116), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n531), .A3(new_n370), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G116), .B(G122), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT93), .A3(new_n370), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n530), .A2(G116), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n370), .B1(new_n539), .B2(KEYINPUT14), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n534), .A2(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n204), .A2(G128), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n203), .A2(G143), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT92), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(G128), .B(G143), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT92), .ZN(new_n547));
  AOI21_X1  g361(.A(G134), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT92), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n544), .A3(new_n221), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n541), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n541), .B(new_n553), .C1(new_n548), .C2(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(KEYINPUT13), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(G134), .C1(KEYINPUT13), .C2(new_n542), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n535), .B(new_n370), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n221), .B1(new_n549), .B2(new_n544), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n528), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n528), .ZN(new_n562));
  INV_X1    g376(.A(new_n560), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n562), .B(new_n563), .C1(new_n552), .C2(new_n554), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n276), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n526), .B1(new_n565), .B2(KEYINPUT95), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(KEYINPUT95), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n568), .B(new_n276), .C1(new_n561), .C2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n570), .B2(new_n526), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n476), .A2(new_n520), .A3(new_n524), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G221), .B1(new_n527), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n250), .A2(G227), .ZN(new_n575));
  XOR2_X1   g389(.A(G110), .B(G140), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n216), .A2(KEYINPUT10), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n446), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n201), .A2(new_n208), .A3(new_n209), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n445), .A2(new_n388), .A3(new_n372), .A4(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT82), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n580), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n408), .A2(new_n237), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT80), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n408), .A2(new_n237), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n417), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n588), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n240), .ZN(new_n595));
  INV_X1    g409(.A(new_n240), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n588), .C1(new_n590), .C2(new_n593), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n578), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT12), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n446), .A2(new_n246), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n600), .A2(new_n582), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n601), .B2(new_n596), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n600), .B2(new_n582), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT12), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(KEYINPUT83), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT83), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n603), .A2(KEYINPUT12), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n599), .B(new_n596), .C1(new_n600), .C2(new_n582), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n597), .A2(new_n605), .A3(new_n609), .A4(new_n578), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n574), .B(new_n276), .C1(new_n598), .C2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n574), .A2(new_n276), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n602), .A2(new_n604), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n597), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n577), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n595), .A2(new_n597), .A3(new_n578), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(G469), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n611), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n468), .A2(new_n572), .A3(new_n573), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n361), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n386), .ZN(G3));
  NAND2_X1  g436(.A1(new_n274), .A2(new_n276), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n279), .A2(new_n281), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n625), .A2(new_n619), .A3(new_n360), .A4(new_n573), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT96), .B1(new_n561), .B2(new_n564), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT96), .B(KEYINPUT33), .C1(new_n561), .C2(new_n564), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n525), .A2(G902), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n631), .A2(new_n632), .B1(new_n525), .B2(new_n565), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n520), .B2(new_n524), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n468), .A2(new_n476), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT34), .B(G104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND2_X1  g452(.A1(new_n468), .A2(new_n476), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n522), .A2(new_n521), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n507), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n276), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n516), .A2(new_n519), .B1(new_n642), .B2(G475), .ZN(new_n643));
  INV_X1    g457(.A(new_n571), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n626), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(new_n620), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n279), .A2(new_n281), .A3(new_n624), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n343), .A2(new_n336), .A3(KEYINPUT97), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT97), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n328), .B2(new_n337), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n653), .A2(new_n655), .B1(KEYINPUT36), .B2(new_n342), .ZN(new_n656));
  INV_X1    g470(.A(new_n653), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT97), .B1(new_n343), .B2(new_n336), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n661), .A2(new_n357), .B1(new_n354), .B2(new_n350), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(new_n573), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n586), .B1(new_n582), .B2(new_n583), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n668), .A2(new_n669), .B1(new_n446), .B2(new_n579), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n592), .A2(new_n591), .A3(new_n417), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT80), .B1(new_n406), .B2(new_n589), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n577), .B1(new_n673), .B2(new_n596), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n674), .A2(new_n595), .B1(new_n615), .B2(new_n577), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n612), .B1(new_n675), .B2(G469), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n667), .B1(new_n676), .B2(new_n611), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n656), .A2(new_n660), .A3(new_n357), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n355), .A2(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n307), .A2(new_n468), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n473), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n471), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n643), .A2(new_n644), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT98), .B(G128), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G30));
  NAND2_X1  g502(.A1(new_n463), .A2(new_n467), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n643), .A2(new_n571), .ZN(new_n692));
  AND4_X1   g506(.A1(new_n362), .A2(new_n691), .A3(new_n662), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n271), .A2(new_n256), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n276), .B1(new_n288), .B2(new_n257), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n282), .A2(new_n283), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n683), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n677), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n698), .B1(new_n700), .B2(KEYINPUT40), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n693), .B(new_n701), .C1(KEYINPUT40), .C2(new_n700), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT100), .B(G143), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G45));
  AOI21_X1  g518(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n517), .A2(KEYINPUT20), .A3(new_n518), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n524), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n633), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n683), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n680), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  OAI21_X1  g525(.A(new_n276), .B1(new_n598), .B2(new_n610), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n573), .A3(new_n611), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n361), .A2(new_n635), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  INV_X1    g531(.A(new_n361), .ZN(new_n718));
  INV_X1    g532(.A(new_n597), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n672), .A2(new_n671), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n596), .B1(new_n720), .B2(new_n588), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n577), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n597), .A2(new_n605), .A3(new_n609), .A4(new_n578), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n574), .B1(new_n724), .B2(new_n276), .ZN(new_n725));
  AOI211_X1 g539(.A(G469), .B(G902), .C1(new_n722), .C2(new_n723), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n726), .A3(new_n667), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n718), .A2(new_n646), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NOR2_X1   g543(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n468), .A3(new_n573), .A4(new_n572), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n307), .A2(new_n679), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT101), .B(G119), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G21));
  NOR2_X1   g549(.A1(G472), .A2(G902), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AND4_X1   g551(.A1(new_n272), .A2(new_n249), .A3(new_n257), .A4(new_n258), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n272), .B1(new_n271), .B2(new_n257), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n287), .A2(new_n289), .A3(new_n293), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n256), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n737), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n359), .A4(new_n475), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n730), .A2(new_n573), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n468), .A2(new_n692), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n530), .ZN(G24));
  NAND3_X1  g563(.A1(new_n707), .A2(new_n708), .A3(new_n683), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n740), .A2(new_n742), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n736), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n624), .A3(new_n679), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n727), .A2(new_n754), .A3(new_n468), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  NAND2_X1  g570(.A1(new_n618), .A2(new_n613), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n573), .B1(new_n726), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n463), .A2(new_n467), .A3(new_n362), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n750), .A2(KEYINPUT42), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n307), .A3(new_n360), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n277), .A2(new_n280), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n296), .A2(new_n299), .A3(new_n276), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n299), .B1(new_n296), .B2(new_n276), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n303), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n283), .B(new_n763), .C1(new_n766), .C2(new_n275), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n677), .A2(new_n360), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n463), .A2(new_n362), .A3(new_n467), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n709), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT42), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(G131), .Z(G33));
  NAND4_X1  g587(.A1(new_n760), .A2(new_n307), .A3(new_n360), .A4(new_n685), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  AOI21_X1  g589(.A(KEYINPUT103), .B1(new_n643), .B2(new_n708), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT43), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n643), .A2(new_n708), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT103), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(KEYINPUT43), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n652), .A3(new_n679), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n616), .A2(new_n617), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n574), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n675), .A2(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n613), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(KEYINPUT102), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT102), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n612), .B1(new_n785), .B2(new_n786), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n726), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n573), .A3(new_n699), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n759), .B(KEYINPUT104), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n782), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n573), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n770), .A2(new_n307), .A3(new_n360), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NAND3_X1  g619(.A1(new_n360), .A2(new_n362), .A3(new_n573), .ZN(new_n806));
  INV_X1    g620(.A(new_n730), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n778), .B(new_n806), .C1(new_n807), .C2(KEYINPUT49), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT105), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(KEYINPUT49), .ZN(new_n810));
  OR4_X1    g624(.A1(new_n691), .A2(new_n809), .A3(new_n697), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n683), .B(KEYINPUT111), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n355), .A2(new_n678), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT112), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n355), .A2(new_n678), .A3(new_n817), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n619), .A2(new_n573), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n747), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n680), .A2(new_n709), .B1(new_n821), .B2(new_n697), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n743), .A2(new_n744), .A3(new_n662), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n634), .A3(new_n683), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n433), .B1(new_n430), .B2(new_n462), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n464), .A2(new_n466), .A3(new_n432), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n362), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n824), .A2(new_n714), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n680), .B2(new_n685), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n813), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n307), .A2(new_n468), .A3(new_n677), .A4(new_n679), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n677), .A2(new_n468), .A3(new_n692), .A4(new_n819), .ZN(new_n832));
  OAI22_X1  g646(.A1(new_n831), .A2(new_n750), .B1(new_n832), .B2(new_n698), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n755), .B1(new_n831), .B2(new_n684), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT113), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n822), .A2(new_n829), .A3(new_n813), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT113), .B1(new_n833), .B2(new_n834), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n626), .A2(new_n639), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n645), .B(KEYINPUT109), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n664), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT106), .B1(new_n643), .B2(new_n633), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT106), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n707), .A2(new_n708), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n468), .A2(new_n846), .A3(new_n476), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT107), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n363), .B(new_n475), .C1(new_n463), .C2(new_n467), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT107), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n846), .A4(new_n848), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n853), .A3(new_n647), .ZN(new_n854));
  INV_X1    g668(.A(new_n621), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n845), .B1(new_n856), .B2(KEYINPUT108), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n731), .A2(new_n732), .B1(new_n746), .B2(new_n747), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n715), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(new_n728), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n707), .A2(new_n644), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n677), .A2(new_n769), .A3(new_n861), .A4(new_n683), .ZN(new_n862));
  INV_X1    g676(.A(new_n732), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(new_n754), .B2(new_n760), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n762), .A2(new_n774), .A3(new_n771), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n626), .B1(new_n849), .B2(KEYINPUT107), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n621), .B1(new_n868), .B2(new_n853), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n857), .A2(new_n860), .A3(new_n867), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n812), .B1(new_n841), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n762), .A2(new_n774), .A3(new_n771), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n728), .A3(new_n859), .A4(new_n864), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n842), .A2(new_n843), .B1(new_n651), .B2(new_n663), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n869), .B2(new_n870), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n856), .A2(KEYINPUT108), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n686), .A2(new_n880), .A3(new_n755), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n822), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n840), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n873), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n840), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n812), .B1(new_n888), .B2(new_n872), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n879), .A2(KEYINPUT53), .A3(new_n840), .A4(new_n836), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n891), .B2(new_n886), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n777), .A2(new_n472), .A3(new_n780), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n777), .A2(KEYINPUT114), .A3(new_n472), .A4(new_n780), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n714), .A2(new_n759), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n359), .A2(new_n471), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n901), .A2(new_n698), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n707), .A2(new_n708), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n902), .A2(new_n823), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n743), .A2(new_n744), .A3(new_n359), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n896), .B2(new_n897), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n691), .A2(new_n362), .A3(new_n714), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(KEYINPUT50), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT50), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n797), .ZN(new_n914));
  INV_X1    g728(.A(new_n802), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n730), .A2(new_n667), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT115), .Z(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n893), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n911), .A2(new_n912), .ZN(new_n920));
  INV_X1    g734(.A(new_n916), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n797), .B(new_n909), .C1(new_n802), .C2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n920), .A2(new_n922), .A3(KEYINPUT51), .A4(new_n906), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n904), .A2(new_n634), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n909), .A2(new_n468), .A3(new_n727), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n924), .A2(new_n469), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n767), .A2(new_n360), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n898), .A2(new_n927), .A3(new_n901), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT48), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n926), .B2(new_n929), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n919), .B(new_n923), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n892), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(G952), .A2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT118), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n811), .B1(new_n934), .B2(new_n936), .ZN(G75));
  NAND2_X1  g751(.A1(new_n873), .A2(new_n885), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(G902), .A3(new_n432), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n423), .B(KEYINPUT119), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT55), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n429), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n939), .B2(new_n940), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n250), .A2(G952), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G51));
  XNOR2_X1  g761(.A(new_n612), .B(KEYINPUT57), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n873), .A2(new_n885), .A3(new_n886), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n886), .B1(new_n873), .B2(new_n885), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n724), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n787), .B(KEYINPUT120), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n938), .A2(G902), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n946), .B1(new_n952), .B2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n938), .A2(G902), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n517), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n517), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n946), .ZN(G60));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n631), .B1(new_n892), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n629), .B2(new_n630), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n949), .B2(new_n950), .ZN(new_n967));
  INV_X1    g781(.A(new_n946), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n965), .A2(new_n969), .ZN(G63));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n873), .B2(new_n885), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n968), .B1(new_n977), .B2(new_n356), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n938), .A2(new_n661), .A3(new_n975), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n938), .A2(new_n975), .ZN(new_n981));
  INV_X1    g795(.A(new_n356), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n977), .A2(new_n661), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(KEYINPUT61), .A3(new_n968), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n985), .ZN(G66));
  INV_X1    g800(.A(G224), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n474), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n857), .A2(new_n860), .A3(new_n871), .ZN(new_n989));
  INV_X1    g803(.A(new_n250), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n941), .B1(G898), .B2(new_n250), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  XOR2_X1   g807(.A(new_n270), .B(KEYINPUT123), .Z(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(new_n509), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(G900), .B(new_n990), .C1(new_n996), .C2(G227), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(G227), .B2(new_n996), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n834), .B(new_n880), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n702), .A3(new_n710), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT124), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n718), .A2(new_n760), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n846), .A2(new_n848), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n699), .B1(new_n843), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n804), .B(new_n798), .C1(new_n1003), .C2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n995), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n999), .A2(new_n710), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n927), .A2(new_n468), .A3(new_n692), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n866), .B1(new_n796), .B2(new_n1013), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n798), .A2(new_n804), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n990), .B1(new_n1015), .B2(new_n996), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n998), .B1(new_n1011), .B2(new_n1016), .ZN(G72));
  INV_X1    g831(.A(new_n694), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1002), .A2(new_n1009), .A3(new_n989), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT126), .ZN(new_n1021));
  XOR2_X1   g835(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  AOI21_X1  g837(.A(new_n1018), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1023), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n1015), .B2(new_n989), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n968), .B1(new_n1026), .B2(new_n301), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1018), .A2(new_n301), .A3(new_n1023), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT127), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n891), .A2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1024), .A2(new_n1027), .A3(new_n1030), .ZN(G57));
endmodule


