

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n554), .A2(n553), .ZN(G160) );
  XOR2_X1 U553 ( .A(KEYINPUT87), .B(n544), .Z(n518) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n660) );
  XNOR2_X1 U555 ( .A(n660), .B(KEYINPUT97), .ZN(n661) );
  XNOR2_X1 U556 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  INV_X1 U558 ( .A(KEYINPUT100), .ZN(n748) );
  NOR2_X1 U559 ( .A1(G2105), .A2(n541), .ZN(n1003) );
  NOR2_X1 U560 ( .A1(G651), .A2(n596), .ZN(n797) );
  NOR2_X1 U561 ( .A1(n545), .A2(n518), .ZN(G164) );
  XOR2_X1 U562 ( .A(G543), .B(KEYINPUT0), .Z(n596) );
  INV_X1 U563 ( .A(G651), .ZN(n527) );
  NOR2_X1 U564 ( .A1(n596), .A2(n527), .ZN(n801) );
  NAND2_X1 U565 ( .A1(G76), .A2(n801), .ZN(n524) );
  XOR2_X1 U566 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n521) );
  NOR2_X1 U567 ( .A1(G543), .A2(G651), .ZN(n519) );
  XNOR2_X1 U568 ( .A(n519), .B(KEYINPUT64), .ZN(n802) );
  NAND2_X1 U569 ( .A1(G89), .A2(n802), .ZN(n520) );
  XNOR2_X1 U570 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U571 ( .A(KEYINPUT74), .B(n522), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U573 ( .A(n525), .B(KEYINPUT5), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n526), .B(KEYINPUT76), .ZN(n535) );
  XNOR2_X1 U575 ( .A(KEYINPUT78), .B(KEYINPUT6), .ZN(n533) );
  NAND2_X1 U576 ( .A1(n797), .A2(G51), .ZN(n531) );
  NOR2_X1 U577 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n528), .Z(n798) );
  NAND2_X1 U579 ( .A1(n798), .A2(G63), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT77), .B(n529), .Z(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U582 ( .A(n533), .B(n532), .Z(n534) );
  NAND2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n536), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n998) );
  NAND2_X1 U586 ( .A1(G114), .A2(n998), .ZN(n538) );
  INV_X1 U587 ( .A(G2104), .ZN(n541) );
  AND2_X1 U588 ( .A1(n541), .A2(G2105), .ZN(n999) );
  NAND2_X1 U589 ( .A1(G126), .A2(n999), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n545) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n539), .Z(n1002) );
  NAND2_X1 U592 ( .A1(n1002), .A2(G138), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n540), .B(KEYINPUT86), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G102), .A2(n1003), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G137), .A2(n1002), .ZN(n547) );
  NAND2_X1 U597 ( .A1(G113), .A2(n998), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n547), .A2(n546), .ZN(n554) );
  NAND2_X1 U599 ( .A1(n999), .A2(G125), .ZN(n548) );
  XNOR2_X1 U600 ( .A(KEYINPUT65), .B(n548), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n1003), .A2(G101), .ZN(n549) );
  XNOR2_X1 U602 ( .A(n549), .B(KEYINPUT23), .ZN(n550) );
  NOR2_X1 U603 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U604 ( .A(KEYINPUT66), .B(n552), .Z(n553) );
  NAND2_X1 U605 ( .A1(G90), .A2(n802), .ZN(n555) );
  XNOR2_X1 U606 ( .A(n555), .B(KEYINPUT70), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G77), .A2(n801), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n557), .A2(n556), .ZN(n559) );
  XOR2_X1 U609 ( .A(KEYINPUT9), .B(KEYINPUT71), .Z(n558) );
  XNOR2_X1 U610 ( .A(n559), .B(n558), .ZN(n563) );
  NAND2_X1 U611 ( .A1(n797), .A2(G52), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G64), .A2(n798), .ZN(n560) );
  AND2_X1 U613 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U614 ( .A1(n563), .A2(n562), .ZN(G301) );
  INV_X1 U615 ( .A(G301), .ZN(G171) );
  NAND2_X1 U616 ( .A1(G75), .A2(n801), .ZN(n565) );
  NAND2_X1 U617 ( .A1(G88), .A2(n802), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U619 ( .A1(G50), .A2(n797), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G62), .A2(n798), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U622 ( .A1(n569), .A2(n568), .ZN(G166) );
  INV_X1 U623 ( .A(G166), .ZN(G303) );
  NAND2_X1 U624 ( .A1(n798), .A2(G65), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G91), .A2(n802), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U627 ( .A1(G78), .A2(n801), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G53), .A2(n797), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U630 ( .A1(n575), .A2(n574), .ZN(G299) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G72), .A2(n801), .ZN(n576) );
  XNOR2_X1 U633 ( .A(n576), .B(KEYINPUT68), .ZN(n579) );
  NAND2_X1 U634 ( .A1(G47), .A2(n797), .ZN(n577) );
  XOR2_X1 U635 ( .A(KEYINPUT69), .B(n577), .Z(n578) );
  NAND2_X1 U636 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G85), .A2(n802), .ZN(n580) );
  XNOR2_X1 U638 ( .A(KEYINPUT67), .B(n580), .ZN(n581) );
  NOR2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U640 ( .A1(n798), .A2(G60), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n584), .A2(n583), .ZN(G290) );
  NAND2_X1 U642 ( .A1(n798), .A2(G61), .ZN(n586) );
  NAND2_X1 U643 ( .A1(G86), .A2(n802), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U645 ( .A(KEYINPUT82), .B(n587), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n801), .A2(G73), .ZN(n588) );
  XOR2_X1 U647 ( .A(KEYINPUT2), .B(n588), .Z(n589) );
  NOR2_X1 U648 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n797), .A2(G48), .ZN(n591) );
  NAND2_X1 U650 ( .A1(n592), .A2(n591), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G49), .A2(n797), .ZN(n594) );
  NAND2_X1 U652 ( .A1(G74), .A2(G651), .ZN(n593) );
  NAND2_X1 U653 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U654 ( .A1(n798), .A2(n595), .ZN(n599) );
  NAND2_X1 U655 ( .A1(G87), .A2(n596), .ZN(n597) );
  XOR2_X1 U656 ( .A(KEYINPUT81), .B(n597), .Z(n598) );
  NAND2_X1 U657 ( .A1(n599), .A2(n598), .ZN(G288) );
  NOR2_X1 U658 ( .A1(G164), .A2(G1384), .ZN(n703) );
  NAND2_X1 U659 ( .A1(G160), .A2(G40), .ZN(n702) );
  INV_X1 U660 ( .A(n702), .ZN(n600) );
  NAND2_X2 U661 ( .A1(n703), .A2(n600), .ZN(n650) );
  NAND2_X1 U662 ( .A1(n650), .A2(G8), .ZN(n601) );
  XOR2_X1 U663 ( .A(KEYINPUT92), .B(n601), .Z(n723) );
  INV_X1 U664 ( .A(n723), .ZN(n718) );
  NOR2_X1 U665 ( .A1(n718), .A2(G1966), .ZN(n676) );
  NOR2_X1 U666 ( .A1(G2084), .A2(n650), .ZN(n675) );
  NOR2_X1 U667 ( .A1(n676), .A2(n675), .ZN(n602) );
  NAND2_X1 U668 ( .A1(G8), .A2(n602), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT30), .ZN(n604) );
  NOR2_X1 U670 ( .A1(G168), .A2(n604), .ZN(n609) );
  INV_X1 U671 ( .A(n650), .ZN(n640) );
  XNOR2_X1 U672 ( .A(G2078), .B(KEYINPUT25), .ZN(n891) );
  NAND2_X1 U673 ( .A1(n640), .A2(n891), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT94), .ZN(n607) );
  OR2_X1 U675 ( .A1(G1961), .A2(n640), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n616) );
  NOR2_X1 U677 ( .A1(G171), .A2(n616), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U679 ( .A(KEYINPUT31), .B(n610), .Z(n673) );
  INV_X1 U680 ( .A(G8), .ZN(n615) );
  NOR2_X1 U681 ( .A1(n718), .A2(G1971), .ZN(n612) );
  NOR2_X1 U682 ( .A1(G2090), .A2(n650), .ZN(n611) );
  NOR2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n613), .A2(G303), .ZN(n614) );
  OR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n667) );
  AND2_X1 U686 ( .A1(n673), .A2(n667), .ZN(n666) );
  AND2_X1 U687 ( .A1(n616), .A2(G171), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n617), .B(KEYINPUT95), .ZN(n664) );
  NAND2_X1 U689 ( .A1(G56), .A2(n798), .ZN(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT14), .B(n618), .Z(n624) );
  NAND2_X1 U691 ( .A1(G81), .A2(n802), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G68), .A2(n801), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U695 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n797), .A2(G43), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n1016) );
  INV_X1 U699 ( .A(G1996), .ZN(n627) );
  NOR2_X1 U700 ( .A1(n650), .A2(n627), .ZN(n628) );
  XOR2_X1 U701 ( .A(n628), .B(KEYINPUT26), .Z(n630) );
  NAND2_X1 U702 ( .A1(n650), .A2(G1341), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n1016), .A2(n631), .ZN(n644) );
  NAND2_X1 U705 ( .A1(n798), .A2(G66), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G92), .A2(n802), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G79), .A2(n801), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G54), .A2(n797), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U712 ( .A(KEYINPUT15), .B(n638), .Z(n639) );
  XNOR2_X1 U713 ( .A(KEYINPUT73), .B(n639), .ZN(n917) );
  NAND2_X1 U714 ( .A1(G1348), .A2(n650), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G2067), .A2(n640), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n917), .A2(n645), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n647) );
  AND2_X1 U719 ( .A1(n917), .A2(n645), .ZN(n646) );
  NOR2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n655) );
  NAND2_X1 U721 ( .A1(n640), .A2(G2072), .ZN(n649) );
  INV_X1 U722 ( .A(KEYINPUT27), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G1956), .A2(n650), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n656) );
  NOR2_X1 U726 ( .A1(G299), .A2(n656), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n653), .B(KEYINPUT96), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U729 ( .A1(G299), .A2(n656), .ZN(n657) );
  XOR2_X1 U730 ( .A(KEYINPUT28), .B(n657), .Z(n658) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(KEYINPUT98), .B(n665), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n666), .A2(n674), .ZN(n671) );
  INV_X1 U735 ( .A(n667), .ZN(n669) );
  AND2_X1 U736 ( .A1(G286), .A2(G8), .ZN(n668) );
  OR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT32), .ZN(n681) );
  AND2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n679) );
  AND2_X1 U741 ( .A1(G8), .A2(n675), .ZN(n677) );
  OR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  OR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n732) );
  NAND2_X1 U745 ( .A1(G166), .A2(G8), .ZN(n682) );
  OR2_X1 U746 ( .A1(G2090), .A2(n682), .ZN(n721) );
  NAND2_X1 U747 ( .A1(G117), .A2(n998), .ZN(n684) );
  NAND2_X1 U748 ( .A1(G129), .A2(n999), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(KEYINPUT89), .ZN(n687) );
  NAND2_X1 U751 ( .A1(G141), .A2(n1002), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n1003), .A2(G105), .ZN(n688) );
  XOR2_X1 U754 ( .A(KEYINPUT38), .B(n688), .Z(n689) );
  NOR2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U756 ( .A(KEYINPUT90), .B(n691), .Z(n995) );
  NAND2_X1 U757 ( .A1(G1996), .A2(n995), .ZN(n699) );
  NAND2_X1 U758 ( .A1(G131), .A2(n1002), .ZN(n693) );
  NAND2_X1 U759 ( .A1(G107), .A2(n998), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U761 ( .A1(G95), .A2(n1003), .ZN(n695) );
  NAND2_X1 U762 ( .A1(G119), .A2(n999), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n990) );
  NAND2_X1 U765 ( .A1(G1991), .A2(n990), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U767 ( .A(KEYINPUT91), .B(n700), .Z(n855) );
  INV_X1 U768 ( .A(n855), .ZN(n701) );
  XOR2_X1 U769 ( .A(G1986), .B(G290), .Z(n916) );
  NAND2_X1 U770 ( .A1(n701), .A2(n916), .ZN(n704) );
  NOR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n760) );
  NAND2_X1 U772 ( .A1(n704), .A2(n760), .ZN(n715) );
  NAND2_X1 U773 ( .A1(n1003), .A2(G104), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n705), .B(KEYINPUT88), .ZN(n707) );
  NAND2_X1 U775 ( .A1(G140), .A2(n1002), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(KEYINPUT34), .B(n708), .ZN(n713) );
  NAND2_X1 U778 ( .A1(G116), .A2(n998), .ZN(n710) );
  NAND2_X1 U779 ( .A1(G128), .A2(n999), .ZN(n709) );
  NAND2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U781 ( .A(KEYINPUT35), .B(n711), .Z(n712) );
  NOR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U783 ( .A(KEYINPUT36), .B(n714), .ZN(n1013) );
  XNOR2_X1 U784 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NOR2_X1 U785 ( .A1(n1013), .A2(n758), .ZN(n849) );
  NAND2_X1 U786 ( .A1(n760), .A2(n849), .ZN(n756) );
  NAND2_X1 U787 ( .A1(n715), .A2(n756), .ZN(n734) );
  NOR2_X1 U788 ( .A1(G1981), .A2(G305), .ZN(n716) );
  XOR2_X1 U789 ( .A(n716), .B(KEYINPUT24), .Z(n717) );
  XNOR2_X1 U790 ( .A(KEYINPUT93), .B(n717), .ZN(n719) );
  INV_X1 U791 ( .A(n718), .ZN(n737) );
  NAND2_X1 U792 ( .A1(n719), .A2(n737), .ZN(n720) );
  OR2_X1 U793 ( .A1(n734), .A2(n720), .ZN(n725) );
  AND2_X1 U794 ( .A1(n721), .A2(n725), .ZN(n722) );
  AND2_X1 U795 ( .A1(n732), .A2(n722), .ZN(n727) );
  OR2_X1 U796 ( .A1(n723), .A2(n734), .ZN(n724) );
  AND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n747) );
  NOR2_X1 U799 ( .A1(G1976), .A2(G288), .ZN(n914) );
  NOR2_X1 U800 ( .A1(G1971), .A2(G303), .ZN(n728) );
  NOR2_X1 U801 ( .A1(n914), .A2(n728), .ZN(n730) );
  INV_X1 U802 ( .A(KEYINPUT33), .ZN(n729) );
  AND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n745) );
  AND2_X1 U805 ( .A1(n914), .A2(KEYINPUT33), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n733), .A2(n737), .ZN(n736) );
  INV_X1 U807 ( .A(n734), .ZN(n735) );
  NAND2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n743) );
  NAND2_X1 U809 ( .A1(G1976), .A2(G288), .ZN(n912) );
  AND2_X1 U810 ( .A1(n737), .A2(n912), .ZN(n738) );
  OR2_X1 U811 ( .A1(KEYINPUT33), .A2(n738), .ZN(n741) );
  XOR2_X1 U812 ( .A(G1981), .B(KEYINPUT99), .Z(n739) );
  XNOR2_X1 U813 ( .A(G305), .B(n739), .ZN(n906) );
  INV_X1 U814 ( .A(n906), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U819 ( .A(n749), .B(n748), .ZN(n763) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n995), .ZN(n750) );
  XOR2_X1 U821 ( .A(KEYINPUT101), .B(n750), .Z(n872) );
  NOR2_X1 U822 ( .A1(G1991), .A2(n990), .ZN(n852) );
  NOR2_X1 U823 ( .A1(G1986), .A2(G290), .ZN(n751) );
  XNOR2_X1 U824 ( .A(KEYINPUT102), .B(n751), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n852), .A2(n752), .ZN(n753) );
  NOR2_X1 U826 ( .A1(n753), .A2(n855), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n872), .A2(n754), .ZN(n755) );
  XNOR2_X1 U828 ( .A(KEYINPUT39), .B(n755), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n1013), .A2(n758), .ZN(n848) );
  NAND2_X1 U831 ( .A1(n759), .A2(n848), .ZN(n761) );
  NAND2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U833 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U834 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U835 ( .A(G2443), .B(G2446), .Z(n766) );
  XNOR2_X1 U836 ( .A(G2427), .B(G2451), .ZN(n765) );
  XNOR2_X1 U837 ( .A(n766), .B(n765), .ZN(n772) );
  XOR2_X1 U838 ( .A(G2430), .B(G2454), .Z(n768) );
  XNOR2_X1 U839 ( .A(G1341), .B(G1348), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n768), .B(n767), .ZN(n770) );
  XOR2_X1 U841 ( .A(G2435), .B(G2438), .Z(n769) );
  XNOR2_X1 U842 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U843 ( .A(n772), .B(n771), .Z(n773) );
  AND2_X1 U844 ( .A1(G14), .A2(n773), .ZN(G401) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U846 ( .A1(G135), .A2(n1002), .ZN(n775) );
  NAND2_X1 U847 ( .A1(G111), .A2(n998), .ZN(n774) );
  NAND2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U849 ( .A1(n999), .A2(G123), .ZN(n776) );
  XOR2_X1 U850 ( .A(KEYINPUT18), .B(n776), .Z(n777) );
  NOR2_X1 U851 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U852 ( .A1(n1003), .A2(G99), .ZN(n779) );
  NAND2_X1 U853 ( .A1(n780), .A2(n779), .ZN(n994) );
  XNOR2_X1 U854 ( .A(G2096), .B(n994), .ZN(n781) );
  OR2_X1 U855 ( .A1(G2100), .A2(n781), .ZN(G156) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  INV_X1 U858 ( .A(G57), .ZN(G237) );
  NAND2_X1 U859 ( .A1(G7), .A2(G661), .ZN(n782) );
  XNOR2_X1 U860 ( .A(n782), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U861 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n784) );
  INV_X1 U862 ( .A(G223), .ZN(n835) );
  NAND2_X1 U863 ( .A1(G567), .A2(n835), .ZN(n783) );
  XNOR2_X1 U864 ( .A(n784), .B(n783), .ZN(G234) );
  INV_X1 U865 ( .A(G860), .ZN(n791) );
  OR2_X1 U866 ( .A1(n1016), .A2(n791), .ZN(G153) );
  NAND2_X1 U867 ( .A1(G868), .A2(G301), .ZN(n786) );
  INV_X1 U868 ( .A(G868), .ZN(n788) );
  NAND2_X1 U869 ( .A1(n917), .A2(n788), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(G284) );
  NOR2_X1 U871 ( .A1(G868), .A2(G299), .ZN(n787) );
  XOR2_X1 U872 ( .A(KEYINPUT79), .B(n787), .Z(n790) );
  NOR2_X1 U873 ( .A1(G286), .A2(n788), .ZN(n789) );
  NOR2_X1 U874 ( .A1(n790), .A2(n789), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n791), .A2(G559), .ZN(n792) );
  INV_X1 U876 ( .A(n917), .ZN(n1019) );
  NAND2_X1 U877 ( .A1(n792), .A2(n1019), .ZN(n793) );
  XNOR2_X1 U878 ( .A(n793), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U879 ( .A1(G868), .A2(n1016), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G868), .A2(n1019), .ZN(n794) );
  NOR2_X1 U881 ( .A1(G559), .A2(n794), .ZN(n795) );
  NOR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(G282) );
  NAND2_X1 U883 ( .A1(G55), .A2(n797), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G67), .A2(n798), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n806) );
  NAND2_X1 U886 ( .A1(G80), .A2(n801), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U889 ( .A1(n806), .A2(n805), .ZN(n817) );
  NAND2_X1 U890 ( .A1(G559), .A2(n1019), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n807), .B(n1016), .ZN(n815) );
  XNOR2_X1 U892 ( .A(KEYINPUT80), .B(n815), .ZN(n808) );
  NOR2_X1 U893 ( .A1(G860), .A2(n808), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n817), .B(n809), .ZN(G145) );
  XNOR2_X1 U895 ( .A(G166), .B(n817), .ZN(n812) );
  XOR2_X1 U896 ( .A(G290), .B(G305), .Z(n810) );
  XNOR2_X1 U897 ( .A(G299), .B(n810), .ZN(n811) );
  XNOR2_X1 U898 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U899 ( .A(KEYINPUT19), .B(n813), .ZN(n814) );
  XNOR2_X1 U900 ( .A(n814), .B(G288), .ZN(n1017) );
  XNOR2_X1 U901 ( .A(n815), .B(n1017), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n816), .A2(G868), .ZN(n819) );
  OR2_X1 U903 ( .A1(n817), .A2(G868), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n821), .ZN(n822) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U909 ( .A1(n823), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U911 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U912 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U913 ( .A1(G108), .A2(n825), .ZN(n963) );
  NAND2_X1 U914 ( .A1(n963), .A2(G567), .ZN(n832) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U917 ( .A1(G218), .A2(n827), .ZN(n828) );
  XOR2_X1 U918 ( .A(KEYINPUT83), .B(n828), .Z(n829) );
  NAND2_X1 U919 ( .A1(G96), .A2(n829), .ZN(n830) );
  XNOR2_X1 U920 ( .A(KEYINPUT84), .B(n830), .ZN(n964) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n964), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n832), .A2(n831), .ZN(n965) );
  NAND2_X1 U923 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U924 ( .A1(n965), .A2(n833), .ZN(n839) );
  NAND2_X1 U925 ( .A1(n839), .A2(G36), .ZN(n834) );
  XOR2_X1 U926 ( .A(KEYINPUT85), .B(n834), .Z(G176) );
  NAND2_X1 U927 ( .A1(n835), .A2(G2106), .ZN(n836) );
  XOR2_X1 U928 ( .A(KEYINPUT103), .B(n836), .Z(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U930 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(G188) );
  NAND2_X1 U934 ( .A1(G124), .A2(n999), .ZN(n840) );
  XOR2_X1 U935 ( .A(KEYINPUT44), .B(n840), .Z(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(KEYINPUT107), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G112), .A2(n998), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U939 ( .A1(G136), .A2(n1002), .ZN(n845) );
  NAND2_X1 U940 ( .A1(G100), .A2(n1003), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U942 ( .A1(n847), .A2(n846), .ZN(G162) );
  INV_X1 U943 ( .A(n848), .ZN(n850) );
  NOR2_X1 U944 ( .A1(n850), .A2(n849), .ZN(n857) );
  XOR2_X1 U945 ( .A(G160), .B(G2084), .Z(n851) );
  NOR2_X1 U946 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U947 ( .A1(n853), .A2(n994), .ZN(n854) );
  NOR2_X1 U948 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U949 ( .A1(n857), .A2(n856), .ZN(n877) );
  NAND2_X1 U950 ( .A1(G139), .A2(n1002), .ZN(n859) );
  NAND2_X1 U951 ( .A1(G103), .A2(n1003), .ZN(n858) );
  NAND2_X1 U952 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U953 ( .A(KEYINPUT108), .B(n860), .ZN(n865) );
  NAND2_X1 U954 ( .A1(G115), .A2(n998), .ZN(n862) );
  NAND2_X1 U955 ( .A1(G127), .A2(n999), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U957 ( .A(KEYINPUT47), .B(n863), .Z(n864) );
  NOR2_X1 U958 ( .A1(n865), .A2(n864), .ZN(n989) );
  XNOR2_X1 U959 ( .A(G2072), .B(n989), .ZN(n868) );
  XNOR2_X1 U960 ( .A(G164), .B(G2078), .ZN(n866) );
  XNOR2_X1 U961 ( .A(n866), .B(KEYINPUT112), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n869), .B(KEYINPUT113), .ZN(n870) );
  XNOR2_X1 U964 ( .A(KEYINPUT50), .B(n870), .ZN(n875) );
  XOR2_X1 U965 ( .A(G2090), .B(G162), .Z(n871) );
  NOR2_X1 U966 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U967 ( .A(KEYINPUT51), .B(n873), .Z(n874) );
  NAND2_X1 U968 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U969 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U970 ( .A(KEYINPUT52), .B(n878), .Z(n879) );
  NOR2_X1 U971 ( .A1(KEYINPUT55), .A2(n879), .ZN(n880) );
  XOR2_X1 U972 ( .A(KEYINPUT114), .B(n880), .Z(n881) );
  NAND2_X1 U973 ( .A1(G29), .A2(n881), .ZN(n961) );
  XNOR2_X1 U974 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n902) );
  XNOR2_X1 U975 ( .A(KEYINPUT115), .B(G2090), .ZN(n882) );
  XNOR2_X1 U976 ( .A(n882), .B(G35), .ZN(n900) );
  XNOR2_X1 U977 ( .A(G1996), .B(G32), .ZN(n884) );
  XNOR2_X1 U978 ( .A(G33), .B(G2072), .ZN(n883) );
  NOR2_X1 U979 ( .A1(n884), .A2(n883), .ZN(n890) );
  XOR2_X1 U980 ( .A(G2067), .B(G26), .Z(n885) );
  NAND2_X1 U981 ( .A1(n885), .A2(G28), .ZN(n888) );
  XNOR2_X1 U982 ( .A(G25), .B(G1991), .ZN(n886) );
  XNOR2_X1 U983 ( .A(KEYINPUT116), .B(n886), .ZN(n887) );
  NOR2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n893) );
  XOR2_X1 U986 ( .A(G27), .B(n891), .Z(n892) );
  NOR2_X1 U987 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U988 ( .A(n894), .B(KEYINPUT117), .Z(n895) );
  XNOR2_X1 U989 ( .A(KEYINPUT53), .B(n895), .ZN(n898) );
  XNOR2_X1 U990 ( .A(G34), .B(G2084), .ZN(n896) );
  XNOR2_X1 U991 ( .A(KEYINPUT54), .B(n896), .ZN(n897) );
  NOR2_X1 U992 ( .A1(n898), .A2(n897), .ZN(n899) );
  NAND2_X1 U993 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n903) );
  OR2_X1 U995 ( .A1(G29), .A2(n903), .ZN(n904) );
  NAND2_X1 U996 ( .A1(G11), .A2(n904), .ZN(n959) );
  XNOR2_X1 U997 ( .A(G16), .B(KEYINPUT56), .ZN(n929) );
  XNOR2_X1 U998 ( .A(G301), .B(G1961), .ZN(n909) );
  XOR2_X1 U999 ( .A(G1966), .B(G168), .Z(n905) );
  NOR2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(KEYINPUT57), .B(n907), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(n909), .A2(n908), .ZN(n927) );
  XNOR2_X1 U1003 ( .A(G1971), .B(G166), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n910), .B(KEYINPUT120), .ZN(n922) );
  XOR2_X1 U1005 ( .A(G1956), .B(G299), .Z(n911) );
  NAND2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n920) );
  XOR2_X1 U1009 ( .A(G1348), .B(n917), .Z(n918) );
  XNOR2_X1 U1010 ( .A(KEYINPUT119), .B(n918), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(n922), .A2(n921), .ZN(n925) );
  XOR2_X1 U1013 ( .A(G1341), .B(n1016), .Z(n923) );
  XNOR2_X1 U1014 ( .A(KEYINPUT121), .B(n923), .ZN(n924) );
  NOR2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1016 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1017 ( .A1(n929), .A2(n928), .ZN(n957) );
  XOR2_X1 U1018 ( .A(G16), .B(KEYINPUT122), .Z(n955) );
  XNOR2_X1 U1019 ( .A(KEYINPUT125), .B(G1966), .ZN(n930) );
  XNOR2_X1 U1020 ( .A(n930), .B(G21), .ZN(n944) );
  XNOR2_X1 U1021 ( .A(G1961), .B(G5), .ZN(n942) );
  XNOR2_X1 U1022 ( .A(G1981), .B(G6), .ZN(n934) );
  XNOR2_X1 U1023 ( .A(KEYINPUT59), .B(G4), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(n931), .B(KEYINPUT123), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(n932), .B(G1348), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1341), .B(G19), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(G1956), .B(G20), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(n939), .B(KEYINPUT60), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(KEYINPUT124), .B(n940), .ZN(n941) );
  NOR2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1035 ( .A(G1971), .B(G22), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(G23), .B(G1976), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1038 ( .A(G1986), .B(KEYINPUT126), .Z(n947) );
  XNOR2_X1 U1039 ( .A(G24), .B(n947), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(KEYINPUT58), .B(n950), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(n953), .B(KEYINPUT61), .ZN(n954) );
  NAND2_X1 U1044 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1045 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1046 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1047 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1048 ( .A(KEYINPUT62), .B(n962), .Z(G311) );
  XNOR2_X1 U1049 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1050 ( .A(G120), .ZN(G236) );
  INV_X1 U1051 ( .A(G96), .ZN(G221) );
  INV_X1 U1052 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(G325) );
  INV_X1 U1054 ( .A(G325), .ZN(G261) );
  INV_X1 U1055 ( .A(n965), .ZN(G319) );
  XOR2_X1 U1056 ( .A(G2100), .B(G2096), .Z(n967) );
  XNOR2_X1 U1057 ( .A(G2072), .B(G2090), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1059 ( .A(G2678), .B(KEYINPUT42), .Z(n969) );
  XNOR2_X1 U1060 ( .A(G2067), .B(KEYINPUT43), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1062 ( .A(n971), .B(n970), .Z(n973) );
  XNOR2_X1 U1063 ( .A(G2084), .B(G2078), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n973), .B(n972), .ZN(G227) );
  XOR2_X1 U1065 ( .A(G2474), .B(KEYINPUT106), .Z(n975) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G1976), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n985) );
  XOR2_X1 U1068 ( .A(G1981), .B(G1986), .Z(n977) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G1991), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n977), .B(n976), .ZN(n981) );
  XOR2_X1 U1071 ( .A(KEYINPUT41), .B(G1971), .Z(n979) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G1956), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n979), .B(n978), .ZN(n980) );
  XOR2_X1 U1074 ( .A(n981), .B(n980), .Z(n983) );
  XNOR2_X1 U1075 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n983), .B(n982), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(n985), .B(n984), .ZN(G229) );
  XOR2_X1 U1078 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n987), .B(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT109), .B(n988), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n994), .B(n993), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n995), .B(G162), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n997), .B(n996), .ZN(n1010) );
  NAND2_X1 U1087 ( .A1(G118), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(G130), .A2(n999), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1008) );
  NAND2_X1 U1090 ( .A1(G142), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(G106), .A2(n1003), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(KEYINPUT45), .B(n1006), .Z(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(n1010), .B(n1009), .Z(n1012) );
  XNOR2_X1 U1096 ( .A(G164), .B(G160), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1012), .B(n1011), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(n1014), .B(n1013), .Z(n1015) );
  NOR2_X1 U1099 ( .A1(G37), .A2(n1015), .ZN(G395) );
  XNOR2_X1 U1100 ( .A(G286), .B(n1016), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(n1018), .B(n1017), .ZN(n1021) );
  XOR2_X1 U1102 ( .A(n1019), .B(G171), .Z(n1020) );
  XNOR2_X1 U1103 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1104 ( .A1(G37), .A2(n1022), .ZN(G397) );
  NOR2_X1 U1105 ( .A1(G227), .A2(G229), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(KEYINPUT49), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(G401), .A2(n1024), .ZN(n1025) );
  AND2_X1 U1108 ( .A1(G319), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1109 ( .A1(G395), .A2(G397), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(G225) );
  INV_X1 U1111 ( .A(G225), .ZN(G308) );
  INV_X1 U1112 ( .A(G108), .ZN(G238) );
endmodule

