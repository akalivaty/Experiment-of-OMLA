//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n469), .B1(new_n474), .B2(new_n468), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n466), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(KEYINPUT70), .B(new_n466), .C1(new_n473), .C2(new_n475), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n471), .A2(new_n470), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n463), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n463), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n487), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT71), .Z(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n470), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n471), .B2(new_n470), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n504), .B(new_n507), .C1(new_n470), .C2(new_n471), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT72), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT73), .Z(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n526), .B1(new_n514), .B2(new_n527), .C1(new_n528), .C2(new_n512), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n512), .A2(new_n531), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n517), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n512), .A2(new_n537), .B1(new_n514), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(new_n512), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n548), .A2(KEYINPUT74), .A3(G91), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  INV_X1    g125(.A(G91), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n512), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n510), .A2(G65), .ZN(new_n554));
  INV_X1    g129(.A(G78), .ZN(new_n555));
  INV_X1    g130(.A(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G299));
  XNOR2_X1  g139(.A(G171), .B(KEYINPUT76), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n548), .A2(G87), .ZN(new_n568));
  INV_X1    g143(.A(new_n514), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n510), .A2(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n517), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI211_X1 g152(.A(KEYINPUT77), .B(new_n517), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n510), .A2(new_n511), .A3(G86), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g156(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n512), .A2(new_n584), .B1(new_n514), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n517), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  AND3_X1   g164(.A1(new_n510), .A2(new_n511), .A3(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n510), .A2(G66), .ZN(new_n592));
  INV_X1    g167(.A(G79), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n556), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n569), .B2(G54), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  MUX2_X1   g172(.A(new_n597), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g173(.A(new_n597), .B(G301), .S(G868), .Z(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g183(.A(KEYINPUT78), .B(KEYINPUT11), .ZN(new_n609));
  XNOR2_X1  g184(.A(G323), .B(new_n609), .ZN(G282));
  XNOR2_X1  g185(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n486), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n490), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n463), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2430), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT81), .Z(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n625), .B2(new_n626), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(G401));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1956), .B(G2474), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1961), .B(G1966), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n652), .A3(new_n653), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n652), .B(new_n653), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n662), .C1(new_n658), .C2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G23), .ZN(new_n672));
  INV_X1    g247(.A(G288), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n673), .B2(new_n671), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT33), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT84), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT32), .B(G1981), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n671), .A2(G6), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n582), .B2(new_n671), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n677), .A2(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n671), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n671), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n677), .B2(new_n678), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n683), .A2(KEYINPUT34), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT34), .B1(new_n683), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n671), .A2(G24), .ZN(new_n691));
  INV_X1    g266(.A(G290), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n671), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n486), .A2(G131), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n490), .A2(G119), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n463), .A2(G107), .ZN(new_n698));
  OAI21_X1  g273(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G25), .B(new_n700), .S(G29), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n689), .A2(new_n690), .A3(new_n695), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT36), .Z(new_n705));
  NAND2_X1  g280(.A1(G162), .A2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G29), .B2(G35), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT29), .Z(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G2090), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(G2090), .ZN(new_n710));
  NOR2_X1   g285(.A1(G5), .A2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT89), .ZN(new_n712));
  INV_X1    g287(.A(G171), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n671), .ZN(new_n714));
  INV_X1    g289(.A(G1961), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT90), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n671), .A2(G4), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n596), .B2(new_n671), .ZN(new_n719));
  INV_X1    g294(.A(G1348), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(new_n463), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n486), .A2(G139), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G33), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G2078), .ZN(new_n734));
  NAND2_X1  g309(.A1(G164), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G27), .B2(G29), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n733), .A2(G2072), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2072), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n732), .A2(new_n738), .B1(new_n715), .B2(new_n714), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n717), .A2(new_n721), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n709), .A2(new_n710), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n730), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n490), .A2(G129), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n486), .A2(G141), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  NAND3_X1  g324(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT87), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(KEYINPUT87), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n743), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n730), .B1(KEYINPUT24), .B2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(KEYINPUT24), .B2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n483), .B2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n756), .A2(new_n757), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n730), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n486), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n490), .A2(G128), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(new_n730), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n671), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n542), .B2(new_n671), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1341), .Z(new_n779));
  XOR2_X1   g354(.A(KEYINPUT31), .B(G11), .Z(new_n780));
  NOR2_X1   g355(.A1(new_n621), .A2(new_n730), .ZN(new_n781));
  INV_X1    g356(.A(G28), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT30), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n782), .B2(KEYINPUT30), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n780), .B(new_n781), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n779), .B(new_n785), .C1(new_n734), .C2(new_n736), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  NOR2_X1   g362(.A1(G168), .A2(new_n671), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n671), .B2(G21), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n776), .B(new_n786), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n787), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT88), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n671), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1956), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n762), .A2(new_n759), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n790), .A2(new_n792), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n705), .A2(new_n742), .A3(new_n766), .A4(new_n798), .ZN(G311));
  INV_X1    g374(.A(G311), .ZN(G150));
  NAND2_X1  g375(.A1(new_n596), .A2(G559), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT92), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT38), .Z(new_n803));
  AND2_X1   g378(.A1(new_n510), .A2(G67), .ZN(new_n804));
  AND2_X1   g379(.A1(G80), .A2(G543), .ZN(new_n805));
  OAI21_X1  g380(.A(G651), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT91), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT91), .ZN(new_n808));
  AOI22_X1  g383(.A1(G93), .A2(new_n548), .B1(new_n569), .B2(G55), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(new_n542), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n803), .B(new_n811), .Z(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(new_n814), .A3(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n817));
  XOR2_X1   g392(.A(new_n816), .B(new_n817), .Z(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n818), .ZN(G145));
  XNOR2_X1  g394(.A(new_n755), .B(new_n773), .ZN(new_n820));
  INV_X1    g395(.A(new_n508), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n507), .B1(new_n474), .B2(new_n504), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n497), .B(new_n501), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n820), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n729), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n490), .A2(G130), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n463), .A2(G118), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G142), .B2(new_n486), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(new_n700), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n613), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT94), .Z(new_n834));
  NOR2_X1   g409(.A1(new_n826), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n483), .B(new_n621), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n495), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n826), .A2(new_n833), .ZN(new_n839));
  AOI21_X1  g414(.A(G37), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n826), .B(new_n834), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT95), .B1(new_n841), .B2(new_n837), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n824), .A2(new_n729), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n824), .A2(new_n729), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n843), .A2(new_n834), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n837), .B1(new_n835), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g423(.A(KEYINPUT40), .B(new_n840), .C1(new_n842), .C2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n841), .A2(KEYINPUT95), .A3(new_n837), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n847), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT40), .B1(new_n853), .B2(new_n840), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n850), .A2(new_n854), .ZN(G395));
  XNOR2_X1  g430(.A(new_n582), .B(G290), .ZN(new_n856));
  XNOR2_X1  g431(.A(G288), .B(G166), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT97), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  INV_X1    g436(.A(new_n858), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(KEYINPUT42), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT98), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n597), .A2(new_n563), .A3(new_n561), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT96), .Z(new_n868));
  NAND2_X1  g443(.A1(G299), .A2(new_n596), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n811), .B(new_n606), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n867), .A2(new_n869), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n865), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n861), .A2(KEYINPUT98), .A3(new_n864), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n865), .A2(new_n879), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n810), .A2(new_n600), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(G295));
  XNOR2_X1  g461(.A(G295), .B(KEYINPUT99), .ZN(G331));
  NOR2_X1   g462(.A1(G168), .A2(G171), .ZN(new_n888));
  INV_X1    g463(.A(G301), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(G168), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n811), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT100), .Z(new_n892));
  OR2_X1    g467(.A1(new_n890), .A2(new_n811), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n892), .A2(new_n878), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n874), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n859), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n859), .B1(new_n895), .B2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n872), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n868), .A2(new_n903), .B1(KEYINPUT41), .B2(new_n878), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n892), .B2(new_n894), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n893), .A2(new_n877), .A3(new_n891), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n860), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n898), .A3(new_n899), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n902), .B1(new_n909), .B2(KEYINPUT43), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT44), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n900), .A2(KEYINPUT43), .A3(new_n901), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n915), .A3(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n917), .B2(KEYINPUT44), .ZN(G397));
  NAND4_X1  g493(.A1(new_n478), .A2(G40), .A3(new_n482), .A4(new_n479), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G164), .B2(G1384), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n755), .A2(G1996), .ZN(new_n923));
  INV_X1    g498(.A(G1996), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n753), .A2(new_n924), .A3(new_n754), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n773), .B(G2067), .Z(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n702), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n700), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n700), .A2(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G290), .B(new_n694), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n922), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n581), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n575), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G1981), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT108), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n943), .A3(G1981), .ZN(new_n944));
  INV_X1    g519(.A(new_n577), .ZN(new_n945));
  INV_X1    g520(.A(G1981), .ZN(new_n946));
  INV_X1    g521(.A(new_n578), .ZN(new_n947));
  INV_X1    g522(.A(new_n581), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n942), .A2(KEYINPUT49), .A3(new_n944), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n949), .A2(new_n944), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(KEYINPUT109), .A3(KEYINPUT49), .A4(new_n942), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n823), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(G8), .B1(new_n919), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n942), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n673), .A2(G1976), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(G8), .C1(new_n919), .C2(new_n957), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n673), .B2(G1976), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(KEYINPUT52), .B2(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n970));
  OAI211_X1 g545(.A(G303), .B(G8), .C1(new_n970), .C2(KEYINPUT55), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT106), .B(KEYINPUT55), .Z(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(G166), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n821), .A2(new_n822), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT45), .B(new_n956), .C1(new_n977), .C2(new_n502), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n921), .A2(KEYINPUT102), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G164), .A2(G1384), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(KEYINPUT45), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n976), .B(new_n919), .C1(new_n979), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n982), .ZN(new_n984));
  INV_X1    g559(.A(new_n919), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT103), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n983), .A2(new_n986), .A3(G1971), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n989), .B(new_n956), .C1(new_n977), .C2(new_n502), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n991), .A2(new_n919), .A3(G2090), .ZN(new_n992));
  OAI21_X1  g567(.A(G8), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n969), .B1(new_n975), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n984), .A2(new_n985), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n976), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n919), .B1(new_n979), .B2(new_n982), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT103), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n686), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT104), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT104), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n1001), .A3(new_n686), .A4(new_n998), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n988), .A2(new_n1003), .A3(new_n990), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n957), .A2(KEYINPUT105), .A3(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n919), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G2090), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1000), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n975), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(G8), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n994), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n919), .A2(G2084), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n921), .A2(new_n978), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n787), .B1(new_n1017), .B2(new_n919), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G286), .A2(G8), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT118), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1021), .B2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1018), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1019), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n1022), .B(KEYINPUT118), .Z(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(KEYINPUT51), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1026), .A3(new_n1031), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1030), .A2(KEYINPUT120), .A3(new_n1031), .A4(new_n1026), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1027), .A2(new_n1034), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1012), .B1(new_n1024), .B2(new_n1039), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1017), .A2(new_n919), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n734), .A2(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1013), .A2(new_n985), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1043), .B1(new_n1048), .B2(new_n715), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n734), .B1(new_n983), .B2(new_n986), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT124), .B1(new_n1055), .B2(new_n889), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1046), .A2(new_n715), .A3(new_n1047), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n480), .A2(KEYINPUT122), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n480), .A2(KEYINPUT122), .ZN(new_n1060));
  AND4_X1   g635(.A1(KEYINPUT53), .A2(new_n482), .A3(G40), .A4(new_n734), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n984), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1057), .B1(new_n1065), .B2(G171), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1058), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1067));
  AOI21_X1  g642(.A(G2078), .B1(new_n996), .B2(new_n998), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT121), .B1(new_n1068), .B2(KEYINPUT53), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(G301), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1056), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1040), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1076), .B2(new_n1049), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n889), .B(new_n1063), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1057), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT123), .ZN(new_n1080));
  OAI211_X1 g655(.A(G301), .B(new_n1064), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1071), .B2(G301), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1057), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  INV_X1    g661(.A(G1956), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n991), .B2(new_n919), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT111), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n1087), .C1(new_n991), .C2(new_n919), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n997), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n553), .A2(new_n563), .A3(KEYINPUT57), .A4(new_n560), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n563), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n563), .A2(new_n1099), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n561), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1095), .A2(new_n1107), .A3(KEYINPUT115), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1089), .A2(new_n1091), .B1(new_n997), .B2(new_n1093), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1106), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1086), .B(new_n1108), .C1(new_n1110), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1109), .A2(KEYINPUT116), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1095), .A2(new_n1107), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1117), .A3(new_n1106), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT61), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n985), .A2(new_n980), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  AOI22_X1  g696(.A1(new_n924), .A2(new_n997), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n542), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1114), .A2(new_n1119), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1114), .A2(new_n1119), .A3(new_n1126), .A4(KEYINPUT117), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1120), .A2(G2067), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1048), .B2(new_n720), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1134), .A2(G1348), .B1(G2067), .B2(new_n1120), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n596), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1129), .A2(new_n1130), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1116), .B1(new_n1132), .B2(new_n597), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1109), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1075), .A2(new_n1085), .A3(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n962), .A2(new_n968), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n999), .A2(KEYINPUT104), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n973), .B(new_n975), .C1(new_n1147), .C2(new_n1002), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1021), .A2(new_n1149), .A3(G8), .A4(G168), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n993), .B2(new_n975), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1010), .B1(new_n1009), .B2(G8), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1030), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1146), .A2(new_n1154), .A3(G168), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT63), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g731(.A(G1976), .B(G288), .C1(new_n955), .C2(new_n961), .ZN(new_n1157));
  INV_X1    g732(.A(new_n949), .ZN(new_n1158));
  OAI211_X1 g733(.A(G8), .B(new_n1120), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n994), .A2(new_n1011), .A3(new_n889), .A4(new_n1055), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1039), .A2(new_n1024), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(KEYINPUT62), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1039), .A2(new_n1164), .A3(new_n1024), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1160), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n935), .B1(new_n1145), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n922), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n924), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT46), .ZN(new_n1170));
  INV_X1    g745(.A(new_n926), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1168), .B1(new_n755), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n930), .B1(new_n927), .B2(new_n1168), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n773), .A2(G2067), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1175), .A2(KEYINPUT125), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT125), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1168), .A3(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n922), .A2(G1986), .A3(G290), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1180), .A2(KEYINPUT48), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(KEYINPUT48), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1181), .B(new_n1182), .C1(new_n933), .C2(new_n922), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1174), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT126), .Z(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT127), .B1(new_n1167), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1055), .A2(new_n889), .ZN(new_n1187));
  AOI211_X1 g762(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1187), .C2(new_n1081), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1083), .B1(new_n1082), .B2(new_n1057), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1074), .B(new_n1040), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1127), .A2(new_n1128), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1191), .A2(new_n1130), .B1(new_n1142), .B2(new_n1109), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1166), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n935), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1185), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1186), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g774(.A1(new_n853), .A2(new_n840), .ZN(new_n1201));
  NOR4_X1   g775(.A1(G401), .A2(new_n461), .A3(G229), .A4(G227), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n1201), .A2(new_n910), .A3(new_n1202), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


