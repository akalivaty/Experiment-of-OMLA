

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U559 ( .A(n634), .B(n633), .ZN(n638) );
  XNOR2_X1 U560 ( .A(n535), .B(n534), .ZN(n536) );
  OR2_X1 U561 ( .A1(n697), .A2(n696), .ZN(n521) );
  AND2_X1 U562 ( .A1(n1002), .A2(n742), .ZN(n522) );
  INV_X1 U563 ( .A(KEYINPUT91), .ZN(n633) );
  INV_X1 U564 ( .A(n660), .ZN(n645) );
  NOR2_X1 U565 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U566 ( .A(n668), .B(KEYINPUT32), .ZN(n676) );
  AND2_X1 U567 ( .A1(n528), .A2(G2104), .ZN(n869) );
  INV_X1 U568 ( .A(KEYINPUT23), .ZN(n534) );
  NOR2_X1 U569 ( .A1(n730), .A2(n522), .ZN(n731) );
  NOR2_X1 U570 ( .A1(n582), .A2(G651), .ZN(n792) );
  AND2_X1 U571 ( .A1(n533), .A2(n532), .ZN(G164) );
  INV_X1 U572 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U573 ( .A1(G102), .A2(n869), .ZN(n525) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n523), .Z(n867) );
  NAND2_X1 U576 ( .A1(G138), .A2(n867), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U578 ( .A(KEYINPUT82), .ZN(n526) );
  XNOR2_X1 U579 ( .A(n527), .B(n526), .ZN(n533) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n528), .ZN(n864) );
  AND2_X1 U581 ( .A1(n864), .A2(G126), .ZN(n531) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n863) );
  NAND2_X1 U583 ( .A1(G114), .A2(n863), .ZN(n529) );
  XNOR2_X1 U584 ( .A(KEYINPUT81), .B(n529), .ZN(n530) );
  NOR2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n864), .A2(G125), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n869), .A2(G101), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U589 ( .A(KEYINPUT64), .B(n538), .ZN(n542) );
  NAND2_X1 U590 ( .A1(G137), .A2(n867), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G113), .A2(n863), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X2 U593 ( .A1(n542), .A2(n541), .ZN(G160) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n582) );
  INV_X1 U595 ( .A(G651), .ZN(n545) );
  NOR2_X1 U596 ( .A1(n582), .A2(n545), .ZN(n784) );
  NAND2_X1 U597 ( .A1(G78), .A2(n784), .ZN(n544) );
  NOR2_X1 U598 ( .A1(G543), .A2(G651), .ZN(n788) );
  NAND2_X1 U599 ( .A1(G91), .A2(n788), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n550) );
  NOR2_X1 U601 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n546), .Z(n547) );
  XNOR2_X1 U603 ( .A(KEYINPUT66), .B(n547), .ZN(n785) );
  NAND2_X1 U604 ( .A1(n785), .A2(G65), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT68), .B(n548), .Z(n549) );
  NOR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n792), .A2(G53), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(G299) );
  NAND2_X1 U609 ( .A1(n792), .A2(G52), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G64), .A2(n785), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U612 ( .A(KEYINPUT67), .B(n555), .Z(n560) );
  NAND2_X1 U613 ( .A1(G77), .A2(n784), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G90), .A2(n788), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U617 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U618 ( .A1(n788), .A2(G89), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G76), .A2(n784), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n564), .B(KEYINPUT5), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n792), .A2(G51), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G63), .A2(n785), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n567), .Z(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U628 ( .A(n570), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G75), .A2(n784), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G88), .A2(n788), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n792), .A2(G50), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G62), .A2(n785), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(n792), .A2(G49), .ZN(n577) );
  XNOR2_X1 U639 ( .A(n577), .B(KEYINPUT76), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT77), .B(n580), .Z(n581) );
  NOR2_X1 U643 ( .A1(n785), .A2(n581), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n582), .A2(G87), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(G288) );
  NAND2_X1 U646 ( .A1(G86), .A2(n788), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G61), .A2(n785), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n784), .A2(G73), .ZN(n587) );
  XOR2_X1 U650 ( .A(KEYINPUT2), .B(n587), .Z(n588) );
  NOR2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n792), .A2(G48), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(G305) );
  NAND2_X1 U654 ( .A1(G85), .A2(n788), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G60), .A2(n785), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U657 ( .A1(G72), .A2(n784), .ZN(n594) );
  XNOR2_X1 U658 ( .A(KEYINPUT65), .B(n594), .ZN(n595) );
  NOR2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U660 ( .A1(n792), .A2(G47), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(G290) );
  NOR2_X1 U662 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n708) );
  INV_X1 U664 ( .A(n708), .ZN(n599) );
  NAND2_X2 U665 ( .A1(n707), .A2(n599), .ZN(n660) );
  NAND2_X1 U666 ( .A1(G8), .A2(n660), .ZN(n693) );
  NAND2_X1 U667 ( .A1(G92), .A2(n788), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G66), .A2(n785), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n606) );
  NAND2_X1 U670 ( .A1(G79), .A2(n784), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G54), .A2(n792), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U673 ( .A(KEYINPUT72), .B(n604), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U675 ( .A(n607), .B(KEYINPUT15), .ZN(n767) );
  NAND2_X1 U676 ( .A1(G1348), .A2(n660), .ZN(n609) );
  NAND2_X1 U677 ( .A1(G2067), .A2(n645), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n609), .A2(n608), .ZN(n626) );
  NOR2_X1 U679 ( .A1(n767), .A2(n626), .ZN(n625) );
  NAND2_X1 U680 ( .A1(n645), .A2(G1996), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT26), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n660), .A2(G1341), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n623) );
  XNOR2_X1 U684 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n788), .A2(G81), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT12), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G68), .A2(n784), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n617), .B(n616), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G56), .A2(n785), .ZN(n618) );
  XOR2_X1 U691 ( .A(KEYINPUT14), .B(n618), .Z(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n792), .A2(G43), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n1011) );
  NOR2_X1 U695 ( .A1(n623), .A2(n1011), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n628) );
  AND2_X1 U697 ( .A1(n767), .A2(n626), .ZN(n627) );
  NOR2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n636) );
  INV_X1 U699 ( .A(KEYINPUT27), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n645), .A2(G2072), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(n632) );
  NAND2_X1 U702 ( .A1(G1956), .A2(n660), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n638), .A2(G299), .ZN(n635) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U706 ( .A(KEYINPUT93), .B(n637), .Z(n642) );
  NAND2_X1 U707 ( .A1(G299), .A2(n638), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n643), .B(KEYINPUT29), .ZN(n650) );
  XOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .Z(n938) );
  NOR2_X1 U712 ( .A1(n938), .A2(n660), .ZN(n644) );
  XOR2_X1 U713 ( .A(KEYINPUT90), .B(n644), .Z(n648) );
  NOR2_X1 U714 ( .A1(n645), .A2(G1961), .ZN(n646) );
  XNOR2_X1 U715 ( .A(KEYINPUT89), .B(n646), .ZN(n647) );
  NAND2_X1 U716 ( .A1(n648), .A2(n647), .ZN(n654) );
  NAND2_X1 U717 ( .A1(G171), .A2(n654), .ZN(n649) );
  NAND2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n659) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n693), .ZN(n672) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n660), .ZN(n669) );
  NOR2_X1 U721 ( .A1(n672), .A2(n669), .ZN(n651) );
  NAND2_X1 U722 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT30), .B(n652), .ZN(n653) );
  NOR2_X1 U724 ( .A1(G168), .A2(n653), .ZN(n656) );
  NOR2_X1 U725 ( .A1(G171), .A2(n654), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT31), .B(n657), .Z(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n670) );
  NAND2_X1 U729 ( .A1(n670), .A2(G286), .ZN(n666) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n693), .ZN(n662) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n660), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT94), .ZN(n664) );
  NAND2_X1 U734 ( .A1(n664), .A2(G303), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U736 ( .A1(n667), .A2(G8), .ZN(n668) );
  NAND2_X1 U737 ( .A1(G8), .A2(n669), .ZN(n674) );
  INV_X1 U738 ( .A(n670), .ZN(n671) );
  NOR2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n688) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n681) );
  NOR2_X1 U743 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n681), .A2(n677), .ZN(n991) );
  NAND2_X1 U745 ( .A1(n688), .A2(n991), .ZN(n678) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NAND2_X1 U747 ( .A1(n678), .A2(n990), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n693), .A2(n679), .ZN(n680) );
  NOR2_X1 U749 ( .A1(KEYINPUT33), .A2(n680), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n681), .A2(KEYINPUT33), .ZN(n682) );
  NOR2_X1 U751 ( .A1(n682), .A2(n693), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(G1981), .B(G305), .Z(n1006) );
  AND2_X1 U754 ( .A1(n685), .A2(n1006), .ZN(n697) );
  NOR2_X1 U755 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U756 ( .A1(G8), .A2(n686), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n689), .A2(n693), .ZN(n695) );
  NOR2_X1 U759 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U760 ( .A(n690), .B(KEYINPUT88), .Z(n691) );
  XNOR2_X1 U761 ( .A(KEYINPUT24), .B(n691), .ZN(n692) );
  OR2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U764 ( .A1(G104), .A2(n869), .ZN(n699) );
  NAND2_X1 U765 ( .A1(G140), .A2(n867), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U767 ( .A(KEYINPUT34), .B(n700), .ZN(n705) );
  NAND2_X1 U768 ( .A1(G116), .A2(n863), .ZN(n702) );
  NAND2_X1 U769 ( .A1(G128), .A2(n864), .ZN(n701) );
  NAND2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U771 ( .A(KEYINPUT35), .B(n703), .Z(n704) );
  NOR2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U773 ( .A(KEYINPUT36), .B(n706), .ZN(n858) );
  XNOR2_X1 U774 ( .A(G2067), .B(KEYINPUT37), .ZN(n739) );
  NOR2_X1 U775 ( .A1(n858), .A2(n739), .ZN(n961) );
  NOR2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n709), .B(KEYINPUT84), .ZN(n742) );
  NAND2_X1 U778 ( .A1(n961), .A2(n742), .ZN(n737) );
  INV_X1 U779 ( .A(n742), .ZN(n727) );
  NAND2_X1 U780 ( .A1(G95), .A2(n869), .ZN(n711) );
  NAND2_X1 U781 ( .A1(G131), .A2(n867), .ZN(n710) );
  NAND2_X1 U782 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U783 ( .A1(G107), .A2(n863), .ZN(n713) );
  NAND2_X1 U784 ( .A1(G119), .A2(n864), .ZN(n712) );
  NAND2_X1 U785 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U786 ( .A1(n715), .A2(n714), .ZN(n857) );
  AND2_X1 U787 ( .A1(n857), .A2(G1991), .ZN(n726) );
  NAND2_X1 U788 ( .A1(n867), .A2(G141), .ZN(n716) );
  XNOR2_X1 U789 ( .A(KEYINPUT86), .B(n716), .ZN(n724) );
  NAND2_X1 U790 ( .A1(G117), .A2(n863), .ZN(n718) );
  NAND2_X1 U791 ( .A1(G129), .A2(n864), .ZN(n717) );
  NAND2_X1 U792 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n869), .A2(G105), .ZN(n719) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n719), .Z(n720) );
  NOR2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U796 ( .A(KEYINPUT85), .B(n722), .Z(n723) );
  NAND2_X1 U797 ( .A1(n724), .A2(n723), .ZN(n851) );
  AND2_X1 U798 ( .A1(G1996), .A2(n851), .ZN(n725) );
  NOR2_X1 U799 ( .A1(n726), .A2(n725), .ZN(n957) );
  NOR2_X1 U800 ( .A1(n727), .A2(n957), .ZN(n734) );
  XNOR2_X1 U801 ( .A(KEYINPUT87), .B(n734), .ZN(n728) );
  NAND2_X1 U802 ( .A1(n737), .A2(n728), .ZN(n730) );
  XOR2_X1 U803 ( .A(G1986), .B(KEYINPUT83), .Z(n729) );
  XNOR2_X1 U804 ( .A(G290), .B(n729), .ZN(n1002) );
  NAND2_X1 U805 ( .A1(n521), .A2(n731), .ZN(n745) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n851), .ZN(n965) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n732) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n857), .ZN(n960) );
  NOR2_X1 U809 ( .A1(n732), .A2(n960), .ZN(n733) );
  NOR2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n965), .A2(n735), .ZN(n736) );
  XNOR2_X1 U812 ( .A(n736), .B(KEYINPUT39), .ZN(n738) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n858), .A2(n739), .ZN(n963) );
  NAND2_X1 U815 ( .A1(n740), .A2(n963), .ZN(n741) );
  XOR2_X1 U816 ( .A(KEYINPUT95), .B(n741), .Z(n743) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U819 ( .A(n746), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U820 ( .A(G2443), .B(G2446), .Z(n748) );
  XNOR2_X1 U821 ( .A(G2451), .B(G2427), .ZN(n747) );
  XNOR2_X1 U822 ( .A(n748), .B(n747), .ZN(n752) );
  XOR2_X1 U823 ( .A(KEYINPUT97), .B(G2454), .Z(n750) );
  XNOR2_X1 U824 ( .A(G2430), .B(G2438), .ZN(n749) );
  XNOR2_X1 U825 ( .A(n750), .B(n749), .ZN(n751) );
  XOR2_X1 U826 ( .A(n752), .B(n751), .Z(n754) );
  XNOR2_X1 U827 ( .A(KEYINPUT98), .B(G2435), .ZN(n753) );
  XNOR2_X1 U828 ( .A(n754), .B(n753), .ZN(n757) );
  XOR2_X1 U829 ( .A(G1341), .B(G1348), .Z(n755) );
  XNOR2_X1 U830 ( .A(KEYINPUT96), .B(n755), .ZN(n756) );
  XOR2_X1 U831 ( .A(n757), .B(n756), .Z(n758) );
  AND2_X1 U832 ( .A1(G14), .A2(n758), .ZN(G401) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  NAND2_X1 U836 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U837 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n761) );
  INV_X1 U839 ( .A(G223), .ZN(n824) );
  NAND2_X1 U840 ( .A1(G567), .A2(n824), .ZN(n760) );
  XNOR2_X1 U841 ( .A(n761), .B(n760), .ZN(G234) );
  INV_X1 U842 ( .A(G860), .ZN(n766) );
  OR2_X1 U843 ( .A1(n1011), .A2(n766), .ZN(G153) );
  INV_X1 U844 ( .A(G171), .ZN(G301) );
  NAND2_X1 U845 ( .A1(G868), .A2(G301), .ZN(n763) );
  INV_X1 U846 ( .A(G868), .ZN(n807) );
  NAND2_X1 U847 ( .A1(n767), .A2(n807), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n763), .A2(n762), .ZN(G284) );
  NOR2_X1 U849 ( .A1(G286), .A2(n807), .ZN(n765) );
  NOR2_X1 U850 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U852 ( .A1(n766), .A2(G559), .ZN(n768) );
  INV_X1 U853 ( .A(n767), .ZN(n998) );
  NAND2_X1 U854 ( .A1(n768), .A2(n998), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n1011), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G868), .A2(n998), .ZN(n770) );
  NOR2_X1 U858 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U860 ( .A1(G99), .A2(n869), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G111), .A2(n863), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n867), .A2(G135), .ZN(n775) );
  XNOR2_X1 U864 ( .A(KEYINPUT73), .B(n775), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n864), .A2(G123), .ZN(n776) );
  XOR2_X1 U866 ( .A(KEYINPUT18), .B(n776), .Z(n777) );
  NOR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U868 ( .A(KEYINPUT74), .B(n779), .Z(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n959) );
  XNOR2_X1 U870 ( .A(n959), .B(G2096), .ZN(n783) );
  INV_X1 U871 ( .A(G2100), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G80), .A2(n784), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G67), .A2(n785), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G93), .A2(n788), .ZN(n789) );
  XNOR2_X1 U877 ( .A(KEYINPUT75), .B(n789), .ZN(n790) );
  NOR2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n792), .A2(G55), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n808) );
  NAND2_X1 U881 ( .A1(n998), .A2(G559), .ZN(n805) );
  XNOR2_X1 U882 ( .A(n1011), .B(n805), .ZN(n795) );
  NOR2_X1 U883 ( .A1(G860), .A2(n795), .ZN(n796) );
  XOR2_X1 U884 ( .A(n808), .B(n796), .Z(G145) );
  XNOR2_X1 U885 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n1011), .B(G166), .ZN(n797) );
  XNOR2_X1 U887 ( .A(n798), .B(n797), .ZN(n799) );
  XNOR2_X1 U888 ( .A(KEYINPUT19), .B(n799), .ZN(n802) );
  XOR2_X1 U889 ( .A(G299), .B(G305), .Z(n800) );
  XNOR2_X1 U890 ( .A(G288), .B(n800), .ZN(n801) );
  XNOR2_X1 U891 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(G290), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(n808), .ZN(n828) );
  XNOR2_X1 U894 ( .A(n828), .B(n805), .ZN(n806) );
  NOR2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n810) );
  NOR2_X1 U896 ( .A1(G868), .A2(n808), .ZN(n809) );
  NOR2_X1 U897 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U900 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U904 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n815) );
  XOR2_X1 U906 ( .A(KEYINPUT22), .B(n815), .Z(n816) );
  NOR2_X1 U907 ( .A1(G218), .A2(n816), .ZN(n817) );
  NAND2_X1 U908 ( .A1(G96), .A2(n817), .ZN(n879) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n879), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT80), .ZN(n822) );
  NAND2_X1 U911 ( .A1(G108), .A2(G120), .ZN(n819) );
  NOR2_X1 U912 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U913 ( .A1(G69), .A2(n820), .ZN(n880) );
  NAND2_X1 U914 ( .A1(G567), .A2(n880), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n881) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n823) );
  NOR2_X1 U917 ( .A1(n881), .A2(n823), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U921 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G120), .B(KEYINPUT99), .ZN(G236) );
  XOR2_X1 U925 ( .A(G96), .B(KEYINPUT100), .Z(G221) );
  XOR2_X1 U926 ( .A(n828), .B(G286), .Z(n830) );
  XNOR2_X1 U927 ( .A(G171), .B(n998), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  NOR2_X1 U929 ( .A1(G37), .A2(n831), .ZN(G397) );
  NAND2_X1 U930 ( .A1(G100), .A2(n869), .ZN(n833) );
  NAND2_X1 U931 ( .A1(G112), .A2(n863), .ZN(n832) );
  NAND2_X1 U932 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n834), .B(KEYINPUT105), .ZN(n836) );
  NAND2_X1 U934 ( .A1(G136), .A2(n867), .ZN(n835) );
  NAND2_X1 U935 ( .A1(n836), .A2(n835), .ZN(n841) );
  XOR2_X1 U936 ( .A(KEYINPUT44), .B(KEYINPUT104), .Z(n838) );
  NAND2_X1 U937 ( .A1(G124), .A2(n864), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(KEYINPUT103), .B(n839), .Z(n840) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G162) );
  NAND2_X1 U941 ( .A1(G103), .A2(n869), .ZN(n843) );
  NAND2_X1 U942 ( .A1(G139), .A2(n867), .ZN(n842) );
  NAND2_X1 U943 ( .A1(n843), .A2(n842), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n864), .A2(G127), .ZN(n844) );
  XNOR2_X1 U945 ( .A(KEYINPUT107), .B(n844), .ZN(n847) );
  NAND2_X1 U946 ( .A1(n863), .A2(G115), .ZN(n845) );
  XOR2_X1 U947 ( .A(KEYINPUT108), .B(n845), .Z(n846) );
  NOR2_X1 U948 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n848), .B(KEYINPUT47), .ZN(n849) );
  NOR2_X1 U950 ( .A1(n850), .A2(n849), .ZN(n974) );
  XNOR2_X1 U951 ( .A(n974), .B(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(G164), .B(G160), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n862) );
  XOR2_X1 U954 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(G162), .B(n856), .ZN(n860) );
  XOR2_X1 U958 ( .A(n858), .B(n857), .Z(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n862), .B(n861), .Z(n877) );
  NAND2_X1 U961 ( .A1(G118), .A2(n863), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G130), .A2(n864), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n874) );
  NAND2_X1 U964 ( .A1(n867), .A2(G142), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT106), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G106), .A2(n869), .ZN(n870) );
  NAND2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n872), .Z(n873) );
  NOR2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U970 ( .A(n959), .B(n875), .ZN(n876) );
  XNOR2_X1 U971 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U972 ( .A1(G37), .A2(n878), .ZN(G395) );
  INV_X1 U974 ( .A(G108), .ZN(G238) );
  INV_X1 U975 ( .A(G69), .ZN(G235) );
  NOR2_X1 U976 ( .A1(n880), .A2(n879), .ZN(G325) );
  INV_X1 U977 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U978 ( .A(KEYINPUT101), .B(n881), .ZN(G319) );
  XOR2_X1 U979 ( .A(G2100), .B(G2096), .Z(n883) );
  XNOR2_X1 U980 ( .A(KEYINPUT42), .B(G2678), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n887) );
  XOR2_X1 U982 ( .A(KEYINPUT43), .B(G2090), .Z(n885) );
  XNOR2_X1 U983 ( .A(G2067), .B(G2072), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U985 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U986 ( .A(G2078), .B(G2084), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(G227) );
  XNOR2_X1 U988 ( .A(G1996), .B(KEYINPUT102), .ZN(n899) );
  XOR2_X1 U989 ( .A(G1976), .B(G1981), .Z(n891) );
  XNOR2_X1 U990 ( .A(G1991), .B(G1966), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U992 ( .A(G1971), .B(G1956), .Z(n893) );
  XNOR2_X1 U993 ( .A(G1986), .B(G1961), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U996 ( .A(G2474), .B(KEYINPUT41), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(G229) );
  XNOR2_X1 U999 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G397), .A2(G395), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n902), .B(KEYINPUT112), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n905), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n906), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1008 ( .A(G1961), .B(G5), .Z(n922) );
  XOR2_X1 U1009 ( .A(G1966), .B(G21), .Z(n907) );
  XNOR2_X1 U1010 ( .A(KEYINPUT125), .B(n907), .ZN(n919) );
  XOR2_X1 U1011 ( .A(KEYINPUT124), .B(G4), .Z(n909) );
  XNOR2_X1 U1012 ( .A(G1348), .B(KEYINPUT59), .ZN(n908) );
  XNOR2_X1 U1013 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1014 ( .A(KEYINPUT123), .B(n910), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(G1341), .B(G19), .ZN(n912) );
  XNOR2_X1 U1016 ( .A(G6), .B(G1981), .ZN(n911) );
  NOR2_X1 U1017 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1018 ( .A1(n914), .A2(n913), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(G20), .B(G1956), .ZN(n915) );
  NOR2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1021 ( .A(KEYINPUT60), .B(n917), .Z(n918) );
  NOR2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(KEYINPUT126), .B(n920), .ZN(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(G1971), .B(G22), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(G23), .B(G1976), .ZN(n923) );
  NOR2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1028 ( .A(G1986), .B(G24), .Z(n925) );
  NAND2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(KEYINPUT58), .B(n927), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(KEYINPUT127), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(KEYINPUT61), .B(n931), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(G16), .A2(n932), .ZN(n956) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n984) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n947) );
  XOR2_X1 U1037 ( .A(G25), .B(G1991), .Z(n933) );
  NAND2_X1 U1038 ( .A1(n933), .A2(G28), .ZN(n944) );
  XOR2_X1 U1039 ( .A(G2067), .B(G26), .Z(n934) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n934), .ZN(n936) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1042 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1043 ( .A(KEYINPUT118), .B(n937), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(G1996), .B(G32), .ZN(n940) );
  XNOR2_X1 U1045 ( .A(n938), .B(G27), .ZN(n939) );
  NOR2_X1 U1046 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1047 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1048 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n945), .ZN(n946) );
  NOR2_X1 U1050 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n948) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n948), .ZN(n949) );
  NAND2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1054 ( .A(n984), .B(n951), .ZN(n953) );
  INV_X1 U1055 ( .A(G29), .ZN(n952) );
  NAND2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n954), .ZN(n955) );
  NOR2_X1 U1058 ( .A1(n956), .A2(n955), .ZN(n988) );
  XNOR2_X1 U1059 ( .A(G160), .B(G2084), .ZN(n958) );
  NAND2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n972) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n970) );
  INV_X1 U1062 ( .A(n961), .ZN(n962) );
  NAND2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n968) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n964) );
  NOR2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(n966), .B(KEYINPUT51), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(KEYINPUT113), .B(n973), .ZN(n982) );
  XOR2_X1 U1071 ( .A(G2072), .B(n974), .Z(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT114), .B(n975), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(G2078), .B(G164), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(KEYINPUT115), .B(n976), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT116), .B(n979), .Z(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT50), .B(n980), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT52), .B(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n986), .A2(G29), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n1018) );
  XOR2_X1 U1083 ( .A(G16), .B(KEYINPUT56), .Z(n1016) );
  XNOR2_X1 U1084 ( .A(G171), .B(G1961), .ZN(n1004) );
  XNOR2_X1 U1085 ( .A(G299), .B(G1956), .ZN(n996) );
  INV_X1 U1086 ( .A(G1971), .ZN(n989) );
  NOR2_X1 U1087 ( .A1(G166), .A2(n989), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1090 ( .A(KEYINPUT119), .B(n994), .ZN(n995) );
  NOR2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1092 ( .A(KEYINPUT120), .B(n997), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n998), .B(G1348), .ZN(n999) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(KEYINPUT121), .B(n1005), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G168), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(n1008), .B(KEYINPUT57), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G1341), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT122), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

