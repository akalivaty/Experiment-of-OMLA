//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  AOI211_X1 g0012(.A(new_n210), .B(new_n212), .C1(G77), .C2(G244), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G1), .B2(G20), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT1), .Z(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR3_X1   g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n220), .A2(new_n217), .A3(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NOR3_X1   g0023(.A1(new_n215), .A2(new_n219), .A3(new_n223), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n226), .B(new_n227), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n245), .B1(G232), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(new_n209), .B2(new_n246), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n248), .B(new_n249), .C1(G107), .C2(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n220), .B(G274), .C1(G41), .C2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G244), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n220), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n251), .B(new_n254), .C1(new_n255), .C2(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(KEYINPUT69), .B(G179), .Z(new_n261));
  OR2_X1    g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G169), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT8), .B(G58), .Z(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n217), .A2(G33), .ZN(new_n269));
  XOR2_X1   g0069(.A(KEYINPUT15), .B(G87), .Z(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n267), .B1(new_n217), .B2(new_n268), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n218), .ZN(new_n274));
  INV_X1    g0074(.A(G13), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n275), .A2(new_n217), .A3(G1), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n272), .A2(new_n274), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n273), .A2(new_n218), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n220), .A2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G77), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n262), .A2(new_n264), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G200), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n246), .A2(G222), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n246), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n250), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(new_n268), .B2(new_n250), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n249), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n252), .B(KEYINPUT66), .ZN(new_n291));
  INV_X1    g0091(.A(new_n259), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(G226), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n283), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(G190), .A3(new_n293), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n203), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n266), .A2(G150), .ZN(new_n298));
  INV_X1    g0098(.A(new_n265), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n297), .B(new_n298), .C1(new_n269), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n274), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n276), .A2(new_n274), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n276), .B2(new_n274), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(G50), .A3(new_n279), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(new_n202), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n295), .A2(new_n296), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(KEYINPUT10), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n294), .B1(new_n311), .B2(new_n308), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n294), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n316), .A2(new_n318), .A3(new_n296), .A4(new_n310), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n261), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n290), .A2(new_n321), .A3(new_n293), .ZN(new_n322));
  AOI21_X1  g0122(.A(G169), .B1(new_n290), .B2(new_n293), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n322), .A2(new_n323), .A3(new_n309), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n260), .A2(G200), .ZN(new_n326));
  INV_X1    g0126(.A(new_n281), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n260), .ZN(new_n329));
  AND4_X1   g0129(.A1(new_n282), .A2(new_n320), .A3(new_n325), .A4(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n303), .A2(new_n265), .A3(new_n279), .A4(new_n305), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n299), .A2(new_n276), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n208), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n266), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n250), .B2(G20), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n342), .B2(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n278), .B1(new_n343), .B2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT73), .B1(new_n243), .B2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT73), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(new_n241), .A3(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(new_n244), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n208), .B1(new_n350), .B2(new_n340), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n351), .B2(new_n338), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n333), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n285), .A2(new_n246), .ZN(new_n354));
  INV_X1    g0154(.A(G226), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n242), .A2(new_n354), .A3(new_n244), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n257), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n291), .ZN(new_n360));
  INV_X1    g0160(.A(G232), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n259), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n328), .A3(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n359), .A2(new_n291), .A3(new_n362), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(G200), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n353), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n353), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n344), .A2(new_n352), .ZN(new_n371));
  INV_X1    g0171(.A(new_n333), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n263), .B1(new_n360), .B2(new_n363), .ZN(new_n374));
  NOR4_X1   g0174(.A1(new_n359), .A2(new_n291), .A3(new_n362), .A4(new_n321), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT18), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n353), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n369), .B(new_n370), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT74), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n266), .A2(G50), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n268), .B2(new_n269), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n217), .A2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n274), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n278), .A2(G68), .A3(new_n279), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n220), .A3(G13), .ZN(new_n391));
  XOR2_X1   g0191(.A(new_n391), .B(KEYINPUT12), .Z(new_n392));
  NOR3_X1   g0192(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n361), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G226), .B2(G1698), .ZN(new_n396));
  INV_X1    g0196(.A(G97), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n245), .B1(new_n241), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n249), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n292), .A2(G238), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n400), .A2(new_n254), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n400), .B2(new_n254), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT13), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n399), .C1(new_n402), .C2(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n328), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n283), .B1(new_n405), .B2(new_n407), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n394), .B(new_n409), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n408), .B2(G169), .ZN(new_n415));
  AOI211_X1 g0215(.A(KEYINPUT14), .B(new_n263), .C1(new_n405), .C2(new_n407), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(G179), .A3(new_n407), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n393), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n330), .A2(new_n382), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G257), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G1698), .ZN(new_n424));
  OR2_X1    g0224(.A1(G250), .A2(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n250), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G294), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n249), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT5), .B(G41), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n220), .A2(G45), .A3(G274), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT82), .ZN(new_n433));
  INV_X1    g0233(.A(G45), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G1), .ZN(new_n435));
  INV_X1    g0235(.A(new_n218), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n430), .A2(new_n435), .B1(new_n436), .B2(new_n256), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n437), .B2(G264), .ZN(new_n438));
  INV_X1    g0238(.A(G41), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT5), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G41), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n435), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G264), .A3(new_n257), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n429), .B(new_n432), .C1(new_n438), .C2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT83), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n437), .A2(new_n433), .A3(G264), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT83), .A3(new_n432), .A4(new_n429), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(G169), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n454));
  INV_X1    g0254(.A(G179), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT84), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n448), .A2(new_n457), .A3(G169), .A4(new_n452), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n220), .A2(G33), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n302), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G20), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n463), .A2(G1), .A3(new_n275), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n461), .A2(new_n462), .B1(KEYINPUT25), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n463), .B(KEYINPUT23), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n242), .A2(new_n244), .A3(new_n217), .A4(G87), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT22), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT81), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n470), .A2(KEYINPUT81), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n467), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n269), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n468), .A2(new_n472), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(new_n477), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT23), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n463), .B(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n250), .A2(new_n217), .A3(new_n471), .A4(G87), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n484), .C1(new_n485), .C2(new_n474), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT24), .B1(new_n486), .B2(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n466), .B1(new_n488), .B2(new_n274), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n465), .A2(KEYINPUT25), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n459), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G190), .B1(new_n448), .B2(new_n452), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n446), .A2(new_n283), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n490), .B(new_n489), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n437), .A2(G257), .B1(new_n431), .B2(new_n430), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n242), .A2(new_n244), .A3(G244), .A4(new_n246), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n246), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT75), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n500), .A2(new_n501), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n506), .A2(KEYINPUT76), .A3(new_n249), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT76), .B1(new_n506), .B2(new_n249), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n249), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G190), .A3(new_n497), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n462), .B1(new_n350), .B2(new_n340), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n266), .A2(G77), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n515), .A2(new_n397), .A3(G107), .ZN(new_n516));
  XNOR2_X1  g0316(.A(G97), .B(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n514), .B1(new_n518), .B2(new_n217), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n274), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n276), .A2(new_n397), .ZN(new_n521));
  INV_X1    g0321(.A(new_n461), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(G97), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n512), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n511), .A2(new_n497), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n263), .A2(new_n525), .B1(new_n520), .B2(new_n523), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n497), .B(new_n321), .C1(new_n507), .C2(new_n508), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n510), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n522), .A2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n276), .A2(new_n478), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n278), .B1(G20), .B2(new_n478), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(new_n241), .B2(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n504), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT20), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT20), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n530), .B(new_n531), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G264), .A2(G1698), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n250), .B(new_n538), .C1(new_n423), .C2(G1698), .ZN(new_n539));
  XOR2_X1   g0339(.A(KEYINPUT79), .B(G303), .Z(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(new_n249), .C1(new_n250), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n437), .A2(G270), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n432), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(G169), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n537), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n543), .A2(new_n328), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n543), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n543), .A2(new_n455), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n537), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n537), .A2(KEYINPUT21), .A3(G169), .A4(new_n543), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n546), .A2(new_n550), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n435), .A2(G274), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT77), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n431), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n257), .B(G250), .C1(G1), .C2(new_n434), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n255), .A2(G1698), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n250), .B(new_n562), .C1(G238), .C2(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G116), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n257), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n250), .A2(new_n217), .A3(G68), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n217), .B1(new_n241), .B2(new_n397), .ZN(new_n569));
  INV_X1    g0369(.A(G87), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n397), .A3(new_n462), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(KEYINPUT19), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n269), .A2(new_n397), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n568), .B(new_n572), .C1(KEYINPUT19), .C2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n274), .B1(new_n276), .B2(new_n271), .ZN(new_n575));
  OAI21_X1  g0375(.A(G200), .B1(new_n561), .B2(new_n565), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n522), .A2(G87), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n567), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n566), .A2(new_n321), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n274), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT78), .B1(new_n461), .B2(new_n271), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n271), .A2(new_n276), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT78), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n302), .A2(new_n583), .A3(new_n460), .A4(new_n270), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n263), .B1(new_n561), .B2(new_n565), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n578), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n529), .A2(new_n554), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n422), .A2(new_n496), .A3(new_n589), .ZN(G372));
  INV_X1    g0390(.A(new_n320), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n353), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT17), .B1(new_n353), .B2(new_n366), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n411), .A2(new_n412), .ZN(new_n596));
  INV_X1    g0396(.A(new_n409), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n393), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n282), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n417), .A2(new_n418), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n394), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n595), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n373), .A2(KEYINPUT18), .A3(new_n377), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n379), .B1(new_n353), .B2(new_n376), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n591), .B1(new_n608), .B2(KEYINPUT87), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n603), .B2(new_n607), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n324), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n492), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n579), .A2(new_n585), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n561), .A2(KEYINPUT85), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n559), .B2(new_n560), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n563), .A2(new_n564), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n617), .A2(new_n619), .B1(new_n257), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n263), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(G200), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n575), .A2(new_n577), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n561), .A2(new_n565), .A3(new_n328), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n495), .A2(new_n528), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n615), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n526), .A2(new_n527), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT26), .B1(new_n588), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n623), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n527), .A2(new_n623), .A3(new_n628), .A4(new_n526), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n613), .B1(new_n459), .B2(new_n491), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n495), .A2(new_n528), .A3(new_n623), .A4(new_n628), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT86), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n631), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n612), .B1(new_n642), .B2(new_n421), .ZN(G369));
  NOR2_X1   g0443(.A1(new_n275), .A2(G20), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n220), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n614), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n459), .A2(new_n491), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n650), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT89), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n491), .A2(new_n650), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n496), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n652), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n492), .A2(new_n650), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n657), .ZN(new_n661));
  INV_X1    g0461(.A(new_n650), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n547), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n613), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n554), .B2(new_n663), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT88), .ZN(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n221), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G1), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n571), .A2(G116), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n216), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n642), .A2(KEYINPUT29), .A3(new_n650), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT92), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n635), .B1(new_n588), .B2(new_n632), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n636), .A2(new_n683), .A3(KEYINPUT26), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT93), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n638), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n495), .A2(new_n528), .A3(new_n628), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n685), .B(new_n623), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n679), .B1(new_n689), .B2(new_n662), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n589), .A2(new_n492), .A3(new_n495), .A4(new_n662), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n496), .A2(KEYINPUT91), .A3(new_n589), .A4(new_n662), .ZN(new_n694));
  INV_X1    g0494(.A(new_n525), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n451), .A2(new_n429), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n551), .A3(new_n696), .A4(new_n566), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT90), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n621), .A2(new_n446), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n543), .A3(new_n509), .A4(new_n321), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n650), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n699), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT31), .B(new_n650), .C1(new_n705), .C2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n693), .A2(new_n694), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n678), .B(new_n690), .C1(G330), .C2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n677), .B1(new_n712), .B2(G1), .ZN(G364));
  AOI21_X1  g0513(.A(new_n218), .B1(G20), .B2(new_n263), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n283), .A2(G179), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G20), .A3(new_n328), .ZN(new_n717));
  INV_X1    g0517(.A(G283), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(G20), .A3(new_n328), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n250), .B1(new_n722), .B2(G329), .ZN(new_n723));
  INV_X1    g0523(.A(G303), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n716), .A2(G20), .A3(G190), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n261), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G190), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G322), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n723), .B1(new_n724), .B2(new_n729), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n731), .A2(new_n328), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT33), .B(G317), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n719), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n732), .A2(new_n283), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n217), .B1(new_n720), .B2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n741), .A2(G326), .B1(G294), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(new_n328), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n740), .B(new_n745), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n729), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G87), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n752), .B(new_n250), .C1(new_n462), .C2(new_n717), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n737), .A2(new_n208), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n742), .A2(new_n397), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n722), .A2(G159), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G58), .A2(new_n733), .B1(new_n748), .B2(G77), .ZN(new_n759));
  INV_X1    g0559(.A(new_n741), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n758), .B(new_n759), .C1(new_n202), .C2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n715), .B1(new_n750), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n714), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n671), .A2(new_n250), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n216), .A2(G45), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n236), .C2(new_n434), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n250), .A2(new_n221), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT94), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G355), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n769), .B(new_n772), .C1(G116), .C2(new_n221), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n762), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n765), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n665), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n674), .B1(G45), .B2(new_n644), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n666), .A2(new_n667), .ZN(new_n779));
  INV_X1    g0579(.A(new_n668), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n778), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n776), .A2(new_n778), .B1(new_n779), .B2(new_n781), .ZN(G396));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n734), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n749), .A2(new_n478), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n729), .A2(new_n462), .B1(new_n397), .B2(new_n742), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n717), .A2(new_n570), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(new_n245), .C1(new_n746), .C2(new_n721), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n737), .A2(KEYINPUT98), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n737), .A2(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n790), .B1(new_n718), .B2(new_n793), .C1(new_n724), .C2(new_n760), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n733), .B1(new_n738), .B2(G150), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n796), .B2(new_n760), .C1(new_n797), .C2(new_n749), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT99), .Z(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n801));
  INV_X1    g0601(.A(new_n717), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G68), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n742), .A2(new_n334), .B1(new_n721), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n751), .B2(G50), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n800), .A2(new_n801), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n794), .B1(new_n807), .B2(new_n245), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n714), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n329), .B1(new_n327), .B2(new_n662), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n282), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n599), .A2(new_n662), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n714), .A2(new_n763), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n813), .A2(new_n763), .B1(new_n268), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n809), .A2(new_n777), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n711), .A2(G330), .ZN(new_n817));
  INV_X1    g0617(.A(new_n813), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n641), .A2(new_n662), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n641), .B2(new_n662), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n817), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n823), .A3(new_n778), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n816), .A2(new_n824), .ZN(G384));
  OAI211_X1 g0625(.A(KEYINPUT31), .B(new_n650), .C1(new_n701), .C2(new_n705), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n693), .A2(new_n694), .A3(new_n708), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n393), .A2(new_n662), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n413), .B2(new_n419), .ZN(new_n829));
  INV_X1    g0629(.A(new_n828), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n602), .A2(new_n598), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n813), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT38), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n208), .B1(new_n340), .B2(new_n341), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n345), .B1(new_n836), .B2(new_n338), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n837), .A3(new_n274), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n372), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(new_n377), .B1(new_n353), .B2(new_n366), .ZN(new_n840));
  INV_X1    g0640(.A(new_n648), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n834), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n371), .A2(new_n372), .B1(new_n376), .B2(new_n648), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n371), .A2(new_n366), .A3(new_n372), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT37), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n842), .B1(new_n594), .B2(new_n606), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n833), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n842), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n381), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n373), .B1(new_n377), .B2(new_n841), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n834), .A3(new_n367), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n839), .A2(new_n377), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n842), .A2(new_n854), .A3(new_n367), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n855), .B2(new_n834), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n851), .A2(new_n856), .A3(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n827), .A2(new_n832), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT40), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n353), .A2(new_n648), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n844), .B2(new_n845), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n381), .A2(new_n863), .B1(new_n853), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n866), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n853), .A2(new_n864), .ZN(new_n869));
  INV_X1    g0669(.A(new_n863), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n594), .B2(new_n606), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT101), .B(new_n868), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n867), .A2(new_n857), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n827), .A2(new_n832), .A3(new_n873), .A4(KEYINPUT40), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n861), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n422), .A2(new_n827), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n875), .B(new_n876), .Z(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(G330), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n819), .A2(new_n812), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n829), .A2(new_n831), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n858), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n602), .A2(new_n650), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n849), .A2(new_n857), .A3(KEYINPUT39), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n606), .A2(new_n841), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n881), .A2(new_n887), .A3(KEYINPUT102), .A4(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n878), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n422), .B1(new_n690), .B2(new_n678), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n612), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n220), .B2(new_n644), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT35), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n217), .B(new_n218), .C1(new_n518), .C2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(G116), .C1(new_n900), .C2(new_n518), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT36), .ZN(new_n903));
  OAI21_X1  g0703(.A(G77), .B1(new_n334), .B2(new_n208), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n904), .A2(new_n216), .B1(G50), .B2(new_n208), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(G1), .A3(new_n275), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT103), .ZN(G367));
  AOI21_X1  g0708(.A(KEYINPUT46), .B1(new_n751), .B2(G116), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n250), .B(new_n909), .C1(G317), .C2(new_n722), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n802), .A2(G97), .B1(new_n743), .B2(G107), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n733), .A2(new_n540), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(G283), .B2(new_n748), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n915), .B1(new_n783), .B2(new_n793), .C1(new_n746), .C2(new_n760), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n717), .A2(new_n268), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n751), .B2(G58), .ZN(new_n918));
  AOI22_X1  g0718(.A1(G143), .A2(new_n741), .B1(new_n733), .B2(G150), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n208), .B2(new_n742), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n918), .B1(new_n797), .B2(new_n793), .C1(new_n920), .C2(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT106), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n245), .B1(new_n722), .B2(G137), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n202), .C2(new_n749), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT47), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n714), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n625), .A2(new_n650), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n623), .A2(new_n628), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n623), .B2(new_n928), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(new_n775), .ZN(new_n931));
  INV_X1    g0731(.A(new_n767), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n766), .B1(new_n221), .B2(new_n271), .C1(new_n232), .C2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n931), .A2(new_n777), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n220), .B1(new_n644), .B2(G45), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n669), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n520), .A2(new_n523), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n528), .B1(new_n939), .B2(new_n662), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n526), .A2(new_n527), .A3(new_n650), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n658), .A2(new_n659), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT44), .B1(new_n660), .B2(new_n942), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n948), .B(new_n943), .C1(new_n658), .C2(new_n659), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n938), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n947), .A2(new_n949), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n944), .B(KEYINPUT45), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n669), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n661), .A2(new_n651), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n658), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(new_n780), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n954), .A3(new_n712), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n712), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n672), .B(KEYINPUT41), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n937), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n938), .A2(new_n942), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n658), .A2(new_n942), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n658), .A2(KEYINPUT42), .A3(new_n942), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n510), .A2(new_n524), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n653), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n650), .B1(new_n971), .B2(new_n632), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n968), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT104), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n972), .B1(new_n966), .B2(new_n967), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT104), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n977), .A3(new_n969), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n976), .A2(new_n969), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n962), .B(new_n963), .C1(new_n979), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n963), .A2(new_n962), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n975), .A2(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n963), .A2(new_n962), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n935), .B1(new_n961), .B2(new_n988), .ZN(G387));
  NAND2_X1  g0789(.A1(new_n957), .A2(new_n937), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n957), .A2(new_n712), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n957), .A2(new_n712), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n672), .A3(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n722), .A2(G326), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G317), .A2(new_n733), .B1(new_n741), .B2(G322), .ZN(new_n996));
  INV_X1    g0796(.A(new_n540), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n996), .B1(new_n997), .B2(new_n749), .C1(new_n793), .C2(new_n746), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT48), .Z(new_n999));
  OAI22_X1  g0799(.A1(new_n729), .A2(new_n783), .B1(new_n718), .B2(new_n742), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT110), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n245), .B1(new_n478), .B2(new_n717), .C1(new_n1002), .C2(KEYINPUT49), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n995), .B(new_n1003), .C1(KEYINPUT49), .C2(new_n1002), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n741), .A2(G159), .B1(G97), .B2(new_n802), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n729), .A2(new_n268), .ZN(new_n1006));
  XOR2_X1   g0806(.A(KEYINPUT108), .B(G150), .Z(new_n1007));
  AOI211_X1 g0807(.A(new_n245), .B(new_n1006), .C1(new_n722), .C2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1005), .B(new_n1008), .C1(new_n208), .C2(new_n749), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n271), .A2(new_n742), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n733), .B2(G50), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT109), .Z(new_n1012));
  AOI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(new_n265), .C2(new_n738), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n714), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n655), .A2(new_n657), .A3(new_n765), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n265), .A2(new_n202), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n675), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n434), .C1(KEYINPUT50), .C2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G68), .B2(G77), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n228), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n767), .B1(new_n1020), .B2(new_n434), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n771), .A2(new_n675), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n221), .A2(G107), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n766), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1014), .A2(new_n777), .A3(new_n1015), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n991), .A2(new_n994), .A3(new_n1026), .ZN(G393));
  NAND2_X1  g0827(.A1(new_n951), .A2(new_n954), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n993), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n672), .A3(new_n958), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n951), .A2(new_n954), .A3(new_n937), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G311), .A2(new_n733), .B1(new_n741), .B2(G317), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  OAI22_X1  g0833(.A1(new_n729), .A2(new_n718), .B1(new_n735), .B2(new_n721), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT111), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1034), .A2(new_n1035), .B1(G107), .B2(new_n802), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n1036), .C1(new_n783), .C2(new_n749), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n250), .B1(new_n743), .B2(G116), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n1035), .B2(new_n1034), .C1(new_n793), .C2(new_n997), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G150), .A2(new_n741), .B1(new_n733), .B2(G159), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n245), .B1(new_n722), .B2(G143), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n268), .B2(new_n742), .C1(new_n749), .C2(new_n299), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n788), .B1(new_n208), .B2(new_n729), .C1(new_n793), .C2(new_n202), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1037), .A2(new_n1039), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n778), .B1(new_n1046), .B2(new_n714), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n766), .B1(new_n397), .B2(new_n221), .C1(new_n239), .C2(new_n932), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n775), .C2(new_n942), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1031), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1030), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT112), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1030), .A2(new_n1050), .A3(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(G390));
  INV_X1    g0855(.A(new_n884), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n689), .A2(new_n662), .A3(new_n811), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1057), .A2(new_n812), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n880), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1056), .B(new_n873), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n884), .B1(new_n879), .B2(new_n880), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n885), .B1(new_n882), .B2(new_n873), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1057), .A2(new_n812), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n884), .B1(new_n1067), .B2(new_n880), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1068), .A2(KEYINPUT113), .A3(new_n873), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n813), .A2(new_n667), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n711), .A2(new_n880), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1062), .A2(new_n1066), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT113), .B1(new_n1068), .B2(new_n873), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1059), .B1(new_n1057), .B2(new_n812), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n873), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1074), .A2(new_n1061), .A3(new_n884), .A4(new_n1075), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1073), .A2(new_n1076), .A3(new_n1065), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n827), .A2(new_n1070), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n1059), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1072), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n422), .A2(G330), .A3(new_n827), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n612), .A2(new_n896), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1078), .A2(new_n1059), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1058), .A2(new_n1071), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n880), .B1(new_n711), .B2(new_n1070), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n879), .B1(new_n1079), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT114), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1082), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1081), .A2(KEYINPUT114), .A3(new_n1091), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n672), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1082), .A2(new_n937), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n245), .B1(new_n722), .B2(G125), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n797), .B2(new_n742), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n751), .A2(new_n1007), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(KEYINPUT53), .B2(new_n1099), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n804), .A2(new_n734), .B1(new_n749), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(G128), .C2(new_n741), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n202), .B2(new_n717), .C1(new_n796), .C2(new_n793), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT115), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n250), .B1(new_n722), .B2(G294), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n749), .B2(new_n397), .C1(new_n718), .C2(new_n760), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n793), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(G107), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n733), .A2(G116), .B1(G77), .B2(new_n743), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT116), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n752), .A3(new_n803), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n715), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n299), .B2(new_n814), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1116), .B(new_n777), .C1(new_n764), .C2(new_n1064), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1095), .A2(new_n1096), .A3(new_n1117), .ZN(G378));
  NAND3_X1  g0918(.A1(new_n861), .A2(G330), .A3(new_n874), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT118), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n320), .B2(new_n325), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(KEYINPUT118), .B(new_n324), .C1(new_n315), .C2(new_n319), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n309), .A2(new_n648), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1119), .B(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n892), .A2(KEYINPUT119), .A3(new_n893), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT119), .B1(new_n892), .B2(new_n893), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT120), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n894), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1133), .B(new_n1140), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1072), .B(new_n1090), .C1(new_n1077), .C2(new_n1080), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1085), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1133), .B(new_n1138), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1144), .A2(new_n1150), .A3(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n672), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1145), .A2(KEYINPUT121), .A3(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1142), .A2(new_n937), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1132), .A2(new_n763), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n814), .A2(new_n202), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n749), .A2(new_n796), .B1(new_n729), .B2(new_n1103), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G150), .B2(new_n743), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G125), .A2(new_n741), .B1(new_n738), .B2(G132), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1161), .C1(new_n1162), .C2(new_n734), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n241), .B1(new_n717), .B2(new_n797), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n1165), .C1(G124), .C2(new_n722), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT117), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1166), .A2(KEYINPUT117), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n462), .A2(new_n734), .B1(new_n760), .B2(new_n478), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n439), .B1(new_n717), .B2(new_n334), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1172), .B(new_n1006), .C1(G283), .C2(new_n722), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n250), .B1(new_n743), .B2(G68), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n749), .C2(new_n271), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1171), .B(new_n1175), .C1(G97), .C2(new_n738), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT58), .Z(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1170), .B(new_n1177), .C1(G50), .C2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n778), .B1(new_n1179), .B2(new_n714), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1157), .A2(new_n1158), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1155), .A2(new_n1183), .ZN(G375));
  NAND3_X1  g0984(.A1(new_n1084), .A2(new_n1089), .A3(new_n1087), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1091), .A2(new_n960), .A3(new_n1185), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n250), .B1(new_n1162), .B2(new_n721), .C1(new_n729), .C2(new_n797), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n717), .A2(new_n334), .B1(new_n742), .B2(new_n202), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n733), .C2(G137), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n748), .A2(G150), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n804), .B2(new_n760), .C1(new_n793), .C2(new_n1103), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n718), .A2(new_n734), .B1(new_n760), .B2(new_n783), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n1010), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n245), .B1(new_n724), .B2(new_n721), .C1(new_n729), .C2(new_n397), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n917), .B(new_n1195), .C1(new_n748), .C2(G107), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(new_n478), .C2(new_n793), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n715), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n778), .B1(new_n208), .B2(new_n814), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT122), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(new_n1059), .C2(new_n763), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1090), .B2(new_n937), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1186), .A2(new_n1202), .ZN(G381));
  NOR2_X1   g1003(.A1(G375), .A2(G378), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G381), .A2(G384), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(G393), .A2(G396), .ZN(new_n1208));
  OR3_X1    g1008(.A1(G390), .A2(G387), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT123), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1206), .A2(new_n1212), .A3(new_n1209), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1211), .A2(new_n1213), .ZN(G407));
  NAND2_X1  g1014(.A1(new_n1204), .A2(new_n649), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G213), .B(new_n1215), .C1(new_n1211), .C2(new_n1213), .ZN(G409));
  INV_X1    g1016(.A(new_n960), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n958), .B2(new_n712), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n987), .B(new_n983), .C1(new_n1218), .C2(new_n937), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1030), .A2(new_n1050), .A3(KEYINPUT112), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT112), .B1(new_n1030), .B2(new_n1050), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n935), .B(new_n1219), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(G387), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT126), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n959), .A2(new_n960), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n936), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n983), .A2(new_n987), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1227), .A2(new_n1228), .B1(new_n934), .B2(new_n927), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(G390), .B2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(G393), .B(G396), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .A4(new_n1231), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1155), .B2(new_n1183), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT125), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1185), .B2(KEYINPUT124), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1185), .A2(new_n1240), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1239), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n672), .B(new_n1091), .C1(new_n1241), .C2(KEYINPUT60), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1202), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G384), .B(new_n1202), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1142), .A2(new_n960), .A3(new_n1144), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1150), .A2(new_n937), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1181), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(G378), .A2(new_n1255), .B1(new_n1256), .B2(G343), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1238), .A2(new_n1252), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1236), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1256), .A2(G343), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(G2897), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1246), .A2(new_n824), .A3(new_n816), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1249), .A3(new_n1262), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1238), .B2(new_n1257), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1257), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT121), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1148), .B(KEYINPUT57), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1182), .B1(new_n1272), .B2(new_n1153), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1251), .B(new_n1269), .C1(new_n1273), .C2(new_n1237), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1235), .B1(new_n1260), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1270), .A2(new_n1271), .A3(new_n1152), .ZN(new_n1278));
  OAI21_X1  g1078(.A(G378), .B1(new_n1278), .B2(new_n1182), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1279), .B2(new_n1269), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1274), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1235), .A2(KEYINPUT61), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1274), .B2(new_n1281), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1238), .A2(new_n1257), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1251), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1282), .A2(new_n1283), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1273), .A2(new_n1237), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1279), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1290), .B1(new_n1291), .B2(new_n1279), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1252), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1235), .B1(new_n1204), .B2(new_n1238), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1251), .A3(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(G402));
endmodule


