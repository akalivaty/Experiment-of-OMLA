//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n459), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g044(.A(new_n469), .B(KEYINPUT65), .Z(G160));
  NAND2_X1  g045(.A1(new_n460), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT66), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n460), .A2(new_n486), .A3(G126), .A4(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n459), .C1(new_n482), .C2(new_n483), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n490), .A2(KEYINPUT67), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n490), .B2(KEYINPUT67), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(G138), .A3(new_n476), .ZN(new_n497));
  INV_X1    g072(.A(G2104), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n488), .A2(new_n492), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n509), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OAI221_X1 g093(.A(new_n506), .B1(new_n507), .B2(new_n514), .C1(new_n518), .C2(new_n508), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  AND2_X1   g095(.A1(new_n505), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  AND3_X1   g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT69), .B(G89), .Z(new_n524));
  OAI221_X1 g099(.A(new_n522), .B1(KEYINPUT7), .B2(new_n523), .C1(new_n514), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(G63), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n508), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n525), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n508), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n505), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(G171));
  NAND4_X1  g115(.A1(new_n509), .A2(new_n511), .A3(G43), .A4(G543), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n514), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(KEYINPUT71), .B(new_n541), .C1(new_n514), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n512), .A2(new_n513), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n545), .A2(new_n546), .B1(G651), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n515), .A2(new_n558), .A3(new_n516), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT73), .B1(new_n512), .B2(new_n513), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(G78), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n535), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n505), .A2(new_n566), .A3(G53), .A4(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n514), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n517), .A2(new_n505), .A3(KEYINPUT72), .A4(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n563), .A2(new_n568), .A3(new_n573), .ZN(G299));
  NAND3_X1  g149(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(G301));
  OAI21_X1  g150(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n517), .A2(new_n505), .A3(G87), .ZN(new_n577));
  AND2_X1   g152(.A1(G49), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT74), .B1(new_n505), .B2(new_n578), .ZN(new_n579));
  AND4_X1   g154(.A1(KEYINPUT74), .A2(new_n509), .A3(new_n511), .A4(new_n578), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n576), .B(new_n577), .C1(new_n579), .C2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n517), .A2(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n508), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n517), .A2(new_n505), .A3(G86), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n505), .A2(G48), .A3(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  NAND3_X1  g164(.A1(new_n505), .A2(G47), .A3(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n517), .A2(new_n505), .A3(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n508), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n514), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n517), .A2(new_n505), .A3(KEYINPUT10), .A4(G92), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n598), .A2(new_n599), .B1(G54), .B2(new_n521), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n559), .B2(new_n560), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT75), .Z(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n600), .A2(KEYINPUT76), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT76), .B1(new_n600), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n595), .B1(new_n594), .B2(new_n608), .ZN(G284));
  XOR2_X1   g184(.A(G284), .B(KEYINPUT77), .Z(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT78), .Z(new_n612));
  AOI21_X1  g187(.A(G868), .B1(G299), .B2(KEYINPUT79), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT79), .B2(G299), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n614), .ZN(G280));
  XOR2_X1   g190(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n607), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n600), .A2(KEYINPUT76), .A3(new_n605), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OR3_X1    g197(.A1(new_n622), .A2(KEYINPUT81), .A3(new_n594), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT81), .B1(new_n622), .B2(new_n594), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n623), .B(new_n624), .C1(G868), .C2(new_n551), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n476), .A2(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT82), .B(G2100), .Z(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n476), .A2(G135), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT83), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n498), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n472), .A2(G123), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n629), .A2(new_n630), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n631), .A2(new_n640), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT86), .Z(new_n665));
  OAI21_X1  g240(.A(new_n663), .B1(new_n662), .B2(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT85), .Z(new_n668));
  INV_X1    g243(.A(new_n663), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n662), .A3(new_n660), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n639), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(G2100), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(G2100), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n679), .B(new_n680), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n678), .B1(KEYINPUT87), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(KEYINPUT87), .B2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NOR2_X1   g270(.A1(G171), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G5), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1961), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(G32), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n472), .A2(G129), .B1(G141), .B2(new_n476), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  NAND3_X1  g279(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n701), .B1(new_n706), .B2(G29), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT27), .B(G1996), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n699), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G2084), .ZN(new_n710));
  NAND2_X1  g285(.A1(G160), .A2(G29), .ZN(new_n711));
  INV_X1    g286(.A(G34), .ZN(new_n712));
  AOI21_X1  g287(.A(G29), .B1(new_n712), .B2(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT24), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n709), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n608), .A2(new_n695), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G4), .B2(new_n695), .ZN(new_n719));
  INV_X1    g294(.A(G1348), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT92), .B(G1341), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n695), .A2(G19), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n551), .B2(new_n695), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n721), .B(new_n722), .C1(new_n723), .C2(new_n726), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n697), .A2(new_n698), .B1(new_n710), .B2(new_n715), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G33), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT94), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n460), .A2(G127), .ZN(new_n731));
  AND2_X1   g306(.A1(G115), .A2(G2104), .ZN(new_n732));
  OAI21_X1  g307(.A(G2105), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n734));
  NAND2_X1  g309(.A1(G103), .A2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n476), .A2(G139), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(new_n700), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n700), .B1(new_n743), .B2(G28), .ZN(new_n745));
  AND2_X1   g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n638), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n707), .A2(new_n708), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n741), .A2(G2072), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n742), .A2(new_n750), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n700), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n700), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2090), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n755), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n476), .A2(G140), .ZN(new_n759));
  NOR2_X1   g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n761));
  INV_X1    g336(.A(G128), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n759), .B1(new_n760), .B2(new_n761), .C1(new_n762), .C2(new_n471), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n700), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n728), .A2(new_n753), .A3(new_n758), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n695), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT23), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n700), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n700), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g353(.A1(G168), .A2(KEYINPUT95), .A3(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(KEYINPUT95), .B1(G168), .B2(G16), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n779), .A2(new_n780), .B1(G16), .B2(G21), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n726), .A2(new_n723), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n769), .A2(new_n778), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n717), .A2(new_n727), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n695), .A2(G6), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n588), .B2(new_n695), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n695), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n695), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G23), .B(G288), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  INV_X1    g374(.A(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT91), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n472), .A2(G119), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT88), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n476), .A2(G131), .ZN(new_n807));
  NOR2_X1   g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G25), .B(new_n810), .S(G29), .Z(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT89), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  MUX2_X1   g391(.A(G24), .B(G290), .S(G16), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1986), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT36), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n821), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n823), .A2(new_n824), .A3(new_n804), .A4(new_n819), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n785), .B1(new_n822), .B2(new_n825), .ZN(G311));
  INV_X1    g401(.A(new_n785), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(G150));
  AOI22_X1  g404(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n508), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n535), .A2(new_n832), .B1(new_n514), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n608), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n550), .A2(G651), .ZN(new_n842));
  INV_X1    g417(.A(new_n546), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n517), .A2(new_n505), .A3(G81), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT71), .B1(new_n844), .B2(new_n541), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g423(.A(KEYINPUT99), .B(new_n842), .C1(new_n843), .C2(new_n845), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n835), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n847), .C1(new_n831), .C2(new_n834), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n841), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT100), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n836), .B1(new_n853), .B2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n838), .B1(new_n855), .B2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(G160), .B(new_n638), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n480), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n476), .A2(G142), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n863), .C1(new_n864), .C2(new_n471), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n628), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n810), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n706), .B(new_n739), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n763), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n493), .A2(new_n495), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n492), .B(new_n502), .C1(new_n489), .C2(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n485), .A2(new_n487), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT101), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n502), .B1(new_n489), .B2(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n488), .A4(new_n492), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n871), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n871), .A2(new_n881), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n869), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n869), .A2(new_n882), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n883), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n888), .A2(new_n885), .A3(new_n868), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n860), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n868), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n859), .A3(new_n886), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT104), .B(G37), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g471(.A1(new_n835), .A2(G868), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n849), .A2(new_n835), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n545), .A2(new_n546), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT99), .B1(new_n899), .B2(new_n842), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n551), .A2(KEYINPUT99), .A3(new_n835), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n621), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n850), .A2(new_n608), .A3(new_n617), .A4(new_n851), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n563), .A2(new_n568), .A3(new_n573), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n600), .A2(new_n605), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT105), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(KEYINPUT105), .A3(new_n906), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n903), .A2(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n600), .A2(new_n605), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(G299), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n910), .A3(new_n918), .A4(new_n915), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n917), .A2(new_n904), .A3(new_n903), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n911), .B1(new_n920), .B2(KEYINPUT106), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n903), .A2(new_n904), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n917), .A4(new_n919), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g503(.A1(G290), .A2(G288), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(G290), .A2(G288), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(KEYINPUT107), .A3(new_n929), .ZN(new_n934));
  XNOR2_X1  g509(.A(G303), .B(new_n588), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n932), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n927), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n935), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n939), .A2(KEYINPUT107), .A3(new_n929), .A4(new_n933), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(KEYINPUT108), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n945), .A3(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n594), .B1(new_n926), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n921), .A2(new_n924), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT109), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n921), .A2(new_n925), .A3(new_n924), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n944), .A2(new_n946), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n897), .B1(new_n954), .B2(KEYINPUT110), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(G295));
  AOI21_X1  g533(.A(KEYINPUT111), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n925), .B1(new_n921), .B2(new_n924), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n926), .A2(new_n960), .A3(new_n947), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n952), .B2(new_n951), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT110), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n897), .ZN(new_n964));
  AND4_X1   g539(.A1(KEYINPUT111), .A2(new_n963), .A3(new_n957), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n959), .A2(new_n965), .ZN(G331));
  NAND2_X1  g541(.A1(new_n917), .A2(new_n919), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n850), .A2(G286), .A3(new_n851), .ZN(new_n968));
  AOI21_X1  g543(.A(G286), .B1(new_n850), .B2(new_n851), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(G171), .ZN(new_n970));
  OAI21_X1  g545(.A(G168), .B1(new_n901), .B2(new_n902), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n850), .A2(G286), .A3(new_n851), .ZN(new_n972));
  AOI21_X1  g547(.A(G301), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(G171), .B1(new_n968), .B2(new_n969), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(G301), .A3(new_n972), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(new_n910), .A3(new_n976), .A4(new_n909), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n943), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n893), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n938), .A2(new_n942), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n970), .A2(new_n973), .A3(new_n916), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n975), .A2(new_n976), .B1(new_n917), .B2(new_n919), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n974), .A2(new_n977), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n980), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n979), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G37), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n978), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n984), .B2(new_n987), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n988), .B2(new_n989), .ZN(new_n997));
  AOI211_X1 g572(.A(KEYINPUT43), .B(new_n992), .C1(new_n984), .C2(new_n987), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT113), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n978), .A2(new_n893), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n986), .B1(new_n985), .B2(new_n980), .ZN(new_n1002));
  AOI211_X1 g577(.A(KEYINPUT112), .B(new_n943), .C1(new_n974), .C2(new_n977), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n995), .B1(new_n1004), .B2(KEYINPUT43), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n993), .A2(new_n989), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n996), .B1(new_n999), .B2(new_n1007), .ZN(G397));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n875), .A2(new_n1009), .A3(new_n879), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n464), .A2(new_n468), .A3(G40), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n706), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2067), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n763), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(KEYINPUT117), .A3(new_n1021), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n810), .A2(new_n814), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n810), .A2(new_n814), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1016), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1024), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(G290), .B2(G1986), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G290), .A2(G1986), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1016), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT61), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n880), .A2(new_n1036), .A3(KEYINPUT45), .A4(new_n1009), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n1009), .A4(new_n879), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT118), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n464), .A2(new_n468), .A3(G40), .ZN(new_n1041));
  INV_X1    g616(.A(new_n492), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(new_n876), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n1043), .B2(new_n488), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1013), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1040), .A2(new_n1041), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n905), .B(KEYINPUT57), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n503), .B2(new_n1009), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT121), .B1(new_n1052), .B2(new_n1015), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n1041), .C1(new_n1044), .C2(new_n1051), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n773), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1049), .A2(new_n1050), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1050), .B1(new_n1049), .B2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1035), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1038), .A2(KEYINPUT118), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1038), .A2(KEYINPUT118), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1041), .B(new_n1047), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1048), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1058), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1050), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1049), .A2(new_n1050), .A3(new_n1058), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(KEYINPUT61), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT58), .B(G1341), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1044), .B2(new_n1041), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1046), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1041), .A2(new_n1017), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT59), .B1(new_n1076), .B2(new_n846), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1046), .B(new_n1074), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1078), .B(new_n551), .C1(new_n1079), .C2(new_n1072), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1044), .A2(new_n1041), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G2067), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n503), .A2(new_n1009), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1015), .B1(new_n1086), .B2(KEYINPUT50), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1087), .A2(new_n1056), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1088), .B2(G1348), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n913), .A2(KEYINPUT60), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1348), .B1(new_n1087), .B2(new_n1056), .ZN(new_n1092));
  NOR4_X1   g667(.A1(new_n1092), .A2(new_n1084), .A3(new_n1082), .A4(new_n1090), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n906), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1092), .A2(new_n1084), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1090), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT126), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(new_n1093), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1061), .A2(new_n1070), .A3(new_n1081), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1099), .A2(new_n906), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1069), .B1(new_n1060), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G166), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT55), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1057), .A2(G2090), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1064), .B2(new_n795), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1113), .B2(new_n1108), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1108), .B1(new_n1044), .B2(new_n1041), .ZN(new_n1116));
  OR2_X1    g691(.A1(G288), .A2(new_n800), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(G288), .B2(new_n800), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1083), .A2(new_n1117), .A3(G8), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n582), .A2(new_n583), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G651), .ZN(new_n1123));
  INV_X1    g698(.A(G1981), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n585), .A4(new_n586), .ZN(new_n1125));
  OAI21_X1  g700(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT49), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1116), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1119), .A2(new_n1121), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT122), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1111), .A2(new_n1108), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1971), .B1(new_n1073), .B2(new_n1041), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1087), .A2(new_n1056), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(G2090), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1134), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1114), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(G301), .B(KEYINPUT54), .ZN(new_n1140));
  INV_X1    g715(.A(G2078), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1041), .A2(KEYINPUT53), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1014), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1064), .B2(G2078), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1144), .B(new_n1146), .C1(G1961), .C2(new_n1088), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n1108), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1966), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1041), .B1(new_n1086), .B2(new_n1013), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1044), .A2(KEYINPUT45), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1087), .A2(new_n710), .A3(new_n1056), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G168), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(G286), .A3(new_n1155), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1150), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1154), .A2(G168), .A3(new_n1155), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT51), .B1(new_n1160), .B2(G8), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1147), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1140), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1073), .A2(new_n1141), .A3(new_n1041), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1165), .A2(new_n1145), .B1(new_n698), .B2(new_n1136), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1044), .A2(KEYINPUT45), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1015), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OR3_X1    g744(.A1(new_n1169), .A2(KEYINPUT127), .A3(G2078), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT127), .B1(new_n1169), .B2(G2078), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(KEYINPUT53), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1164), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1139), .A2(new_n1163), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1107), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1154), .A2(G286), .A3(new_n1155), .ZN(new_n1178));
  AOI21_X1  g753(.A(G286), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1149), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1160), .A2(G8), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1180), .B(KEYINPUT62), .C1(KEYINPUT51), .C2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1172), .B(new_n1146), .C1(G1961), .C2(new_n1088), .ZN(new_n1183));
  AND4_X1   g758(.A1(G171), .A2(new_n1177), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1139), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G288), .A2(G1976), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1131), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1125), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1116), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1131), .A2(new_n1121), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT119), .B1(new_n1190), .B2(new_n1118), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1119), .A2(new_n1192), .A3(new_n1121), .A4(new_n1131), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1189), .B1(new_n1138), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(KEYINPUT120), .B(new_n1189), .C1(new_n1138), .C2(new_n1195), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1184), .A2(new_n1185), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1175), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1157), .A2(new_n1108), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1114), .A2(new_n1133), .A3(new_n1138), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n1204));
  XNOR2_X1  g779(.A(KEYINPUT123), .B(KEYINPUT63), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1204), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1110), .A2(KEYINPUT125), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1194), .A2(KEYINPUT63), .A3(new_n1202), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1206), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1034), .B1(new_n1201), .B2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1014), .A2(G1996), .A3(new_n1015), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n1216), .A2(KEYINPUT46), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(KEYINPUT46), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1020), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1016), .B1(new_n706), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT47), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1223), .B1(G2067), .B2(new_n763), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1016), .ZN(new_n1225));
  NOR4_X1   g800(.A1(new_n1014), .A2(G1986), .A3(G290), .A4(new_n1015), .ZN(new_n1226));
  XOR2_X1   g801(.A(new_n1226), .B(KEYINPUT48), .Z(new_n1227));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n1029), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1222), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1215), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g805(.A1(new_n674), .A2(G319), .A3(new_n658), .A4(new_n675), .ZN(new_n1232));
  AOI211_X1 g806(.A(G229), .B(new_n1232), .C1(new_n890), .C2(new_n894), .ZN(new_n1233));
  AND2_X1   g807(.A1(new_n1233), .A2(new_n994), .ZN(G308));
  NAND2_X1  g808(.A1(new_n1233), .A2(new_n994), .ZN(G225));
endmodule


