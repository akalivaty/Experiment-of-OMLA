//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT72), .B(G902), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  OAI211_X1 g005(.A(G134), .B(new_n190), .C1(new_n191), .C2(KEYINPUT65), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n193), .B(KEYINPUT11), .C1(new_n194), .C2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n190), .A2(KEYINPUT67), .A3(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G137), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n198), .A2(KEYINPUT67), .B1(KEYINPUT65), .B2(new_n191), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n199), .A3(new_n202), .A4(new_n197), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT76), .A3(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n211), .A2(new_n205), .A3(KEYINPUT76), .A4(G104), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n208), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n205), .A3(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT77), .B1(new_n205), .B2(G104), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n209), .A2(G107), .ZN(new_n217));
  OAI211_X1 g031(.A(G101), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(KEYINPUT64), .A3(G143), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT64), .B1(new_n224), .B2(G143), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n221), .B(new_n223), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(G143), .B2(new_n224), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n231), .B2(new_n222), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n219), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n213), .A2(new_n218), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n222), .B2(new_n231), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n227), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n204), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(KEYINPUT12), .B(new_n204), .C1(new_n234), .C2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n207), .A2(new_n210), .A3(new_n212), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n220), .B2(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n224), .A2(KEYINPUT64), .A3(G143), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n248), .A2(new_n249), .B1(new_n220), .B2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n221), .B2(new_n228), .ZN(new_n253));
  OR2_X1    g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n250), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n244), .A2(new_n256), .A3(G101), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n246), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n204), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n238), .B2(KEYINPUT10), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n231), .A2(new_n222), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n227), .B1(new_n250), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n219), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(KEYINPUT78), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n260), .A2(new_n261), .A3(new_n263), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G110), .B(G140), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G227), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n243), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n263), .A2(new_n258), .A3(new_n259), .A4(new_n268), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n204), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n273), .B1(new_n277), .B2(new_n269), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n187), .B(new_n189), .C1(new_n275), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n243), .A2(new_n269), .ZN(new_n280));
  INV_X1    g094(.A(new_n273), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n277), .A2(new_n269), .A3(new_n273), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(G469), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(G469), .A2(G902), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G221), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT9), .B(G234), .Z(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  XOR2_X1   g107(.A(G116), .B(G119), .Z(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT2), .B(G113), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n246), .A2(new_n296), .A3(new_n257), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G116), .ZN(new_n301));
  OAI211_X1 g115(.A(G113), .B(new_n301), .C1(new_n294), .C2(new_n299), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n219), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G110), .B(G122), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n297), .A2(new_n303), .A3(new_n305), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(KEYINPUT6), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G224), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G953), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n227), .A2(new_n232), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n255), .A2(new_n312), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(KEYINPUT79), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n229), .A2(new_n251), .A3(new_n254), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n236), .B2(new_n251), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n311), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(KEYINPUT79), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n319), .ZN(new_n323));
  INV_X1    g137(.A(new_n311), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n313), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n304), .A2(new_n327), .A3(new_n306), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n309), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G210), .B1(G237), .B2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(new_n313), .A3(KEYINPUT80), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT81), .B(KEYINPUT7), .Z(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n324), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n332), .B(new_n334), .C1(KEYINPUT80), .C2(new_n313), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n305), .B(KEYINPUT8), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n302), .A2(new_n298), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n337), .A2(new_n235), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n235), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n340), .A3(new_n308), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT7), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n325), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n289), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n329), .A2(new_n331), .A3(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n335), .A2(new_n340), .A3(new_n308), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n325), .A2(new_n342), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n309), .A2(new_n326), .A3(new_n328), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n330), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n293), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n292), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n312), .A2(KEYINPUT16), .A3(G140), .ZN(new_n354));
  XNOR2_X1  g168(.A(G125), .B(G140), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G146), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT19), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g173(.A1(G125), .A2(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(G125), .A2(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT19), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n224), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n202), .ZN(new_n365));
  OR2_X1    g179(.A1(KEYINPUT69), .A2(G237), .ZN(new_n366));
  NAND2_X1  g180(.A1(KEYINPUT69), .A2(G237), .ZN(new_n367));
  AOI21_X1  g181(.A(G953), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G143), .B1(new_n368), .B2(G214), .ZN(new_n369));
  AND2_X1   g183(.A1(KEYINPUT69), .A2(G237), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT69), .A2(G237), .ZN(new_n371));
  OAI211_X1 g185(.A(G214), .B(new_n271), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n220), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n365), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n220), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT69), .B(G237), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n376), .A2(G143), .A3(G214), .A4(new_n271), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n377), .A3(new_n202), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n364), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT18), .ZN(new_n382));
  INV_X1    g196(.A(G131), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT82), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n375), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n375), .B2(new_n377), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n355), .B(new_n224), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n381), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n384), .B1(new_n369), .B2(new_n373), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n375), .A2(new_n377), .A3(new_n385), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n391), .A2(new_n381), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n380), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n209), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n389), .A3(new_n392), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n379), .B1(new_n402), .B2(new_n393), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT84), .B1(new_n403), .B2(new_n398), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n356), .A2(G146), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n356), .A2(G146), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n202), .B1(new_n375), .B2(new_n377), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n405), .B(new_n406), .C1(KEYINPUT17), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n374), .A2(new_n409), .A3(new_n378), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n374), .A2(KEYINPUT85), .A3(new_n409), .A4(new_n378), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n402), .A2(new_n393), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n398), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n400), .A2(new_n404), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n417), .A2(KEYINPUT86), .A3(new_n420), .A4(new_n422), .ZN(new_n425));
  INV_X1    g239(.A(new_n416), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n398), .B1(new_n414), .B2(new_n415), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n289), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n424), .A2(new_n425), .B1(G475), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT87), .B1(new_n220), .B2(G128), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n222), .A3(G143), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n220), .A2(G128), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n194), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT88), .ZN(new_n442));
  AOI21_X1  g256(.A(G134), .B1(new_n442), .B2(new_n437), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n430), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G116), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n445), .A2(G122), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(KEYINPUT90), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n447), .B2(new_n446), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n445), .A2(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n451), .A2(KEYINPUT90), .B1(new_n446), .B2(new_n447), .ZN(new_n452));
  OAI21_X1  g266(.A(G107), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(KEYINPUT91), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n194), .B1(new_n438), .B2(new_n439), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n442), .A2(G134), .A3(new_n437), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT89), .A3(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n446), .A2(new_n450), .A3(G107), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n453), .B2(KEYINPUT91), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n444), .A2(new_n454), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n436), .B(KEYINPUT13), .Z(new_n461));
  INV_X1    g275(.A(new_n434), .ZN(new_n462));
  OAI21_X1  g276(.A(G134), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n446), .A2(new_n450), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n205), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n455), .B(new_n463), .C1(new_n465), .C2(new_n458), .ZN(new_n466));
  INV_X1    g280(.A(new_n288), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT73), .B(G217), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n467), .A2(G953), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n460), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n460), .B2(new_n466), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT92), .B(new_n189), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G478), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT15), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n460), .A2(new_n466), .ZN(new_n478));
  INV_X1    g292(.A(new_n470), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n471), .ZN(new_n481));
  INV_X1    g295(.A(new_n476), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(KEYINPUT92), .A3(new_n189), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n271), .A2(G952), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(G234), .B2(G237), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT21), .B(G898), .Z(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT93), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(G234), .A2(G237), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n188), .A2(G953), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n485), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n477), .A2(new_n483), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n353), .B1(new_n429), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n428), .A2(G475), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n419), .A2(new_n420), .B1(new_n417), .B2(new_n422), .ZN(new_n498));
  INV_X1    g312(.A(new_n425), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n500), .A2(KEYINPUT94), .A3(new_n494), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n352), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT95), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n429), .A2(new_n353), .A3(new_n495), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT94), .B1(new_n500), .B2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT95), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n352), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(G101), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n368), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT70), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n317), .B1(new_n201), .B2(new_n203), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT68), .B1(new_n194), .B2(G137), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n190), .A3(G134), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n517), .A3(new_n198), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G131), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n233), .A2(new_n203), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n296), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT28), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  NOR4_X1   g338(.A1(new_n514), .A2(new_n520), .A3(new_n524), .A4(new_n296), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n296), .B1(new_n514), .B2(new_n520), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n513), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n204), .A2(new_n255), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n233), .A2(new_n203), .A3(new_n519), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n514), .A2(new_n520), .A3(KEYINPUT30), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n296), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n522), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n512), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n514), .A2(new_n520), .A3(new_n296), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n529), .A3(new_n531), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT30), .B1(new_n514), .B2(new_n520), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(new_n296), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT31), .A3(new_n512), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n528), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G472), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT32), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n523), .ZN(new_n549));
  INV_X1    g363(.A(new_n525), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n527), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n513), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT31), .B1(new_n543), .B2(new_n512), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n522), .B1(new_n540), .B2(new_n541), .ZN(new_n555));
  INV_X1    g369(.A(new_n512), .ZN(new_n556));
  NOR4_X1   g370(.A1(new_n555), .A2(new_n537), .A3(new_n539), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT32), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n546), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n535), .A2(new_n561), .A3(new_n527), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT71), .B(new_n296), .C1(new_n514), .C2(new_n520), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT28), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n564), .A2(KEYINPUT29), .A3(new_n512), .A4(new_n549), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT29), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n551), .B2(new_n552), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n543), .A2(new_n512), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n189), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n548), .A2(new_n560), .B1(G472), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT25), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n300), .A2(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n222), .A2(G119), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(G119), .B2(new_n222), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n300), .A2(KEYINPUT23), .A3(G128), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G110), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n575), .B(new_n580), .C1(new_n406), .C2(new_n405), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n355), .A2(new_n224), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(G110), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n582), .B(new_n357), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n581), .A2(KEYINPUT75), .A3(new_n585), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT74), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n271), .A2(G221), .A3(G234), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n586), .A3(new_n587), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n571), .B1(new_n597), .B2(new_n189), .ZN(new_n598));
  AOI211_X1 g412(.A(KEYINPUT25), .B(new_n188), .C1(new_n594), .C2(new_n596), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n469), .B1(new_n189), .B2(G234), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(G902), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n600), .A2(new_n601), .B1(new_n602), .B2(new_n597), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n570), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n503), .A2(new_n508), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n472), .B2(new_n473), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n480), .A2(KEYINPUT98), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(KEYINPUT33), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n188), .A2(new_n475), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n481), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n481), .A2(new_n189), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n475), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n500), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n351), .A2(KEYINPUT96), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n331), .B1(new_n329), .B2(new_n344), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n348), .A2(new_n330), .A3(new_n349), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n293), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n619), .A2(new_n626), .A3(new_n492), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n545), .B2(new_n188), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n547), .B2(new_n545), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n629), .A2(new_n604), .A3(new_n292), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n631), .B(new_n633), .ZN(G6));
  AOI21_X1  g448(.A(new_n624), .B1(new_n623), .B2(new_n293), .ZN(new_n635));
  INV_X1    g449(.A(new_n293), .ZN(new_n636));
  AOI211_X1 g450(.A(KEYINPUT96), .B(new_n636), .C1(new_n621), .C2(new_n622), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n492), .B1(new_n477), .B2(new_n483), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n423), .A2(new_n420), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n417), .A2(KEYINPUT20), .A3(new_n422), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n640), .A2(new_n497), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n638), .A2(KEYINPUT100), .A3(new_n639), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n620), .A2(new_n642), .A3(new_n625), .A4(new_n639), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n630), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(new_n629), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n586), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n655), .A2(new_n602), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n600), .B2(new_n601), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n503), .A2(new_n508), .A3(new_n653), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT37), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(G12));
  NAND2_X1  g475(.A1(new_n569), .A2(G472), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n545), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n559), .B1(new_n558), .B2(new_n546), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n286), .A2(new_n291), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n620), .A4(new_n625), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n485), .B(KEYINPUT104), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT103), .B(G900), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n491), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n640), .A2(new_n497), .A3(new_n641), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n477), .A2(new_n483), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n658), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT105), .B1(new_n667), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n570), .A2(new_n292), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n477), .A2(new_n483), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n673), .A2(new_n680), .A3(new_n657), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n678), .A2(new_n679), .A3(new_n638), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XOR2_X1   g498(.A(new_n672), .B(KEYINPUT39), .Z(new_n685));
  NOR2_X1   g499(.A1(new_n292), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT40), .Z(new_n687));
  OR2_X1    g501(.A1(new_n623), .A2(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n623), .A2(KEYINPUT106), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(KEYINPUT38), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT38), .B1(new_n688), .B2(new_n689), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n293), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n552), .A2(new_n563), .A3(new_n562), .ZN(new_n694));
  INV_X1    g508(.A(new_n536), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n289), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n663), .B2(new_n664), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n675), .A3(new_n500), .A4(new_n657), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n693), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n700), .B1(new_n693), .B2(new_n699), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n687), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n220), .ZN(G45));
  NAND4_X1  g519(.A1(new_n500), .A2(new_n618), .A3(new_n658), .A4(new_n672), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n667), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n224), .ZN(G48));
  AND2_X1   g522(.A1(new_n277), .A2(new_n269), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n274), .B1(new_n709), .B2(new_n273), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n189), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n291), .A3(new_n279), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n570), .A2(new_n713), .A3(new_n604), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n627), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT108), .B(KEYINPUT109), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  INV_X1    g533(.A(new_n713), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n665), .A3(new_n603), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n643), .B2(new_n646), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n445), .ZN(G18));
  NOR3_X1   g537(.A1(new_n626), .A2(new_n713), .A3(new_n657), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n506), .A2(new_n724), .A3(new_n665), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND2_X1  g540(.A1(new_n638), .A2(new_n639), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n564), .A2(new_n549), .ZN(new_n728));
  OAI22_X1  g542(.A1(new_n728), .A2(new_n513), .B1(new_n554), .B2(new_n557), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n546), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n558), .A2(new_n189), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n731), .B1(new_n732), .B2(G472), .ZN(new_n733));
  INV_X1    g547(.A(G472), .ZN(new_n734));
  AOI211_X1 g548(.A(KEYINPUT110), .B(new_n734), .C1(new_n558), .C2(new_n189), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n603), .B(new_n730), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n628), .A2(KEYINPUT110), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n732), .A2(new_n731), .A3(G472), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(KEYINPUT111), .A3(new_n603), .A4(new_n730), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n727), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n429), .A2(new_n713), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  AND3_X1   g560(.A1(new_n500), .A2(new_n618), .A3(new_n672), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n739), .A2(new_n740), .B1(new_n546), .B2(new_n729), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n720), .A2(new_n638), .A3(new_n658), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n724), .A2(new_n752), .A3(new_n747), .A4(new_n748), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n282), .A2(KEYINPUT113), .A3(G469), .A4(new_n283), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n279), .A2(new_n759), .A3(new_n285), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n284), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n290), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n621), .A2(new_n293), .A3(new_n622), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n665), .A3(new_n603), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n756), .A2(new_n757), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n500), .A2(new_n618), .A3(new_n672), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n758), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n570), .A2(new_n604), .A3(new_n764), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n500), .A2(new_n618), .A3(new_n672), .A4(new_n767), .ZN(new_n771));
  INV_X1    g585(.A(new_n758), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n763), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n383), .ZN(G33));
  NAND4_X1  g589(.A1(new_n770), .A2(new_n675), .A3(new_n674), .A4(new_n763), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  AND2_X1   g591(.A1(new_n615), .A2(new_n617), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n500), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n778), .B2(new_n500), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n629), .A3(new_n658), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n282), .A2(new_n283), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n282), .A2(KEYINPUT45), .A3(new_n283), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(G469), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n285), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(KEYINPUT46), .A3(new_n285), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n279), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n291), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n685), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n784), .A2(new_n785), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n786), .A2(new_n765), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT115), .B(G137), .Z(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(G39));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n796), .B2(new_n291), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n806), .A2(new_n603), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n672), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n619), .A2(new_n665), .A3(new_n811), .A4(new_n764), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(KEYINPUT117), .A3(new_n812), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NOR3_X1   g632(.A1(new_n692), .A2(new_n604), .A3(new_n698), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n712), .A2(new_n279), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n293), .B1(new_n820), .B2(KEYINPUT49), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(KEYINPUT49), .B2(new_n820), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n291), .A3(new_n779), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n698), .A2(new_n604), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n713), .A2(new_n764), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n485), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT122), .A4(new_n485), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n429), .A3(new_n778), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n669), .B1(new_n780), .B2(new_n782), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n658), .A3(new_n748), .A4(new_n825), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n636), .B(new_n720), .C1(new_n690), .C2(new_n691), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n738), .A2(new_n742), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n831), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n833), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n831), .A2(new_n837), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(new_n765), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n712), .A2(new_n290), .A3(new_n279), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n806), .B2(new_n809), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT123), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n847), .A2(KEYINPUT123), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n839), .B(new_n840), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n765), .A3(new_n844), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT51), .B1(new_n854), .B2(KEYINPUT120), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n833), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n844), .A2(new_n638), .A3(new_n720), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n500), .A2(new_n618), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n828), .A2(new_n860), .A3(new_n829), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n831), .A2(new_n605), .A3(new_n825), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n484), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n858), .A2(new_n859), .A3(new_n861), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n722), .B1(new_n743), .B2(new_n744), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n769), .A2(new_n773), .A3(new_n776), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n725), .A2(new_n715), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n747), .A2(new_n748), .A3(new_n763), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n675), .B(KEYINPUT119), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n666), .A2(new_n872), .A3(new_n665), .A4(new_n674), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n658), .B(new_n765), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n619), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n876), .B(new_n878), .C1(new_n500), .C2(new_n872), .ZN(new_n879));
  INV_X1    g693(.A(new_n351), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n493), .A3(new_n880), .A4(new_n630), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n659), .A2(new_n881), .A3(new_n606), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n707), .B1(new_n677), .B2(new_n682), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n626), .A2(new_n429), .A3(new_n680), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n658), .A2(new_n811), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n698), .A3(new_n763), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n754), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n754), .A2(new_n884), .A3(KEYINPUT52), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n883), .A2(new_n892), .A3(KEYINPUT53), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT53), .B1(new_n883), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n867), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n893), .A2(new_n894), .A3(new_n867), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n866), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n823), .B1(new_n897), .B2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n271), .A2(G952), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n309), .A2(new_n328), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n326), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT55), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n188), .B(new_n331), .C1(new_n893), .C2(new_n894), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n188), .B1(new_n893), .B2(new_n894), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT125), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n188), .C1(new_n893), .C2(new_n894), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n331), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT126), .B(KEYINPUT56), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n903), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n900), .B(new_n907), .C1(new_n912), .C2(new_n914), .ZN(G51));
  XOR2_X1   g729(.A(new_n285), .B(KEYINPUT57), .Z(new_n916));
  NAND3_X1  g730(.A1(new_n896), .A2(new_n895), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n710), .ZN(new_n918));
  INV_X1    g732(.A(new_n791), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n909), .A2(new_n919), .A3(new_n911), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n900), .B1(new_n918), .B2(new_n920), .ZN(G54));
  AND2_X1   g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n909), .A2(new_n911), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n417), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n900), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n909), .A2(new_n417), .A3(new_n911), .A4(new_n922), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT59), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n896), .A2(new_n895), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n611), .A2(new_n614), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n896), .A2(new_n932), .A3(new_n895), .A4(new_n930), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(new_n926), .A3(new_n935), .ZN(G63));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n893), .A2(new_n894), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n655), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n926), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n597), .B1(new_n938), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n938), .A2(new_n940), .ZN(new_n945));
  INV_X1    g759(.A(new_n597), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n926), .A4(new_n941), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n488), .B2(new_n310), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n868), .A2(new_n870), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n882), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n901), .B1(G898), .B2(new_n271), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  AND2_X1   g769(.A1(new_n359), .A2(new_n362), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n542), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(G900), .B1(new_n957), .B2(G227), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n271), .B(new_n958), .C1(G227), .C2(new_n957), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n786), .A2(new_n765), .A3(new_n799), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n885), .A2(new_n605), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n798), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n754), .A2(new_n884), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n817), .A3(new_n869), .A4(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n957), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n704), .B2(new_n964), .ZN(new_n971));
  INV_X1    g785(.A(new_n703), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n701), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT62), .B(new_n965), .C1(new_n973), .C2(new_n687), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n879), .A2(new_n686), .A3(new_n770), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n817), .A2(new_n800), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n967), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n959), .B1(new_n969), .B2(new_n980), .ZN(G72));
  OR2_X1    g795(.A1(new_n695), .A2(new_n568), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n512), .B1(new_n975), .B2(new_n979), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n966), .A2(new_n556), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n984), .A3(new_n952), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n938), .A2(new_n982), .A3(new_n987), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n900), .A3(new_n989), .ZN(G57));
endmodule


