//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G8gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  OR2_X1    g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G57gat), .B(G64gat), .Z(new_n214));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n209), .B2(new_n211), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n210), .A2(KEYINPUT89), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT90), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n216), .A2(KEYINPUT90), .A3(new_n217), .A4(new_n218), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n213), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n207), .B1(new_n223), .B2(KEYINPUT21), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G231gat), .A2(G233gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G155gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n228), .B(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n223), .A2(KEYINPUT21), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT91), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT92), .B(G183gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n236), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OR3_X1    g039(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n242), .B1(G29gat), .B2(G36gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT15), .ZN(new_n244));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245));
  OR3_X1    g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n245), .A2(new_n244), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n244), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT17), .ZN(new_n251));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252));
  INV_X1    g051(.A(G85gat), .ZN(new_n253));
  INV_X1    g052(.A(G92gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(KEYINPUT8), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT7), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n253), .B2(new_n254), .ZN(new_n257));
  NAND3_X1  g056(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G99gat), .B(G106gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT94), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n255), .A2(new_n260), .A3(new_n257), .A4(new_n258), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n264), .A2(new_n263), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT93), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT41), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n267), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G190gat), .B(G218gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n272), .A2(KEYINPUT41), .ZN(new_n278));
  XNOR2_X1  g077(.A(G134gat), .B(G162gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT95), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n278), .B(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n277), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n240), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT82), .B(G22gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT71), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n289));
  OR2_X1    g088(.A1(G197gat), .A2(G204gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n288), .B(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n286), .B1(new_n293), .B2(KEYINPUT29), .ZN(new_n294));
  INV_X1    g093(.A(G155gat), .ZN(new_n295));
  INV_X1    g094(.A(G162gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT74), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G155gat), .B2(G162gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n297), .A2(new_n299), .B1(G155gat), .B2(G162gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G141gat), .B(G148gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(KEYINPUT2), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(KEYINPUT75), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G141gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n296), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(KEYINPUT2), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n302), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n302), .A2(new_n313), .A3(new_n286), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n293), .B1(KEYINPUT29), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n317), .B1(new_n315), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n285), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT84), .ZN(new_n324));
  INV_X1    g123(.A(new_n322), .ZN(new_n325));
  INV_X1    g124(.A(new_n285), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n320), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT83), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n320), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n285), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n325), .A2(new_n332), .A3(new_n320), .A4(new_n326), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n324), .A2(new_n328), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335));
  INV_X1    g134(.A(G50gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n329), .A2(G22gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n339), .A3(new_n327), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT66), .Z(new_n348));
  OAI211_X1 g147(.A(new_n345), .B(new_n346), .C1(new_n348), .C2(KEYINPUT26), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT27), .B(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT68), .B1(new_n352), .B2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n353), .A2(new_n354), .B1(G183gat), .B2(G190gat), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n352), .A2(KEYINPUT68), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n356), .A2(new_n353), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n349), .B(new_n355), .C1(new_n357), .C2(new_n354), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n347), .B1(KEYINPUT65), .B2(new_n359), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n359), .A2(KEYINPUT65), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n360), .A2(new_n361), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT23), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(KEYINPUT25), .ZN(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n366), .A2(new_n351), .A3(KEYINPUT24), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n351), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n362), .B(new_n371), .C1(new_n348), .C2(new_n359), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n365), .A2(new_n371), .B1(new_n372), .B2(KEYINPUT25), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G120gat), .ZN(new_n377));
  INV_X1    g176(.A(G120gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G113gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT69), .B1(new_n377), .B2(new_n379), .ZN(new_n381));
  AND2_X1   g180(.A1(G127gat), .A2(G134gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(G127gat), .A2(G134gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G113gat), .B(G120gat), .Z(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n375), .C1(KEYINPUT69), .C2(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n386), .A2(new_n388), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n358), .A2(new_n391), .A3(new_n373), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n394), .B(KEYINPUT64), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n395), .A3(new_n392), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT32), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT32), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n400), .A3(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G15gat), .B(G43gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n398), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT33), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n403), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n399), .A2(new_n411), .A3(new_n401), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n410), .B1(new_n404), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n344), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417));
  INV_X1    g216(.A(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT72), .B(G8gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n374), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n358), .B2(new_n373), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n293), .ZN(new_n427));
  INV_X1    g226(.A(new_n293), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n424), .B(new_n428), .C1(new_n423), .C2(new_n425), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n422), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT73), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n422), .A3(new_n429), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT35), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT77), .ZN(new_n437));
  AND4_X1   g236(.A1(KEYINPUT4), .A2(new_n389), .A3(new_n302), .A4(new_n313), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n307), .A2(G141gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n305), .A2(G148gat), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT75), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT75), .B1(new_n439), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n443), .A2(new_n312), .B1(new_n444), .B2(new_n300), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT4), .B1(new_n445), .B2(new_n389), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n437), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n286), .B1(new_n302), .B2(new_n313), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n318), .A2(new_n448), .A3(new_n389), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT76), .Z(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n445), .A2(KEYINPUT77), .A3(new_n454), .A4(new_n389), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n447), .A2(new_n450), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n391), .B2(new_n314), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n445), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n449), .B1(new_n460), .B2(new_n437), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n453), .A4(new_n455), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n391), .A2(new_n314), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n389), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n452), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n452), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT5), .B(new_n468), .C1(new_n470), .C2(new_n460), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G85gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT0), .B(G57gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n476), .A3(new_n471), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n435), .A2(new_n436), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n416), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n478), .A2(KEYINPUT79), .A3(new_n479), .A4(new_n482), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n481), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n491), .A2(new_n492), .A3(new_n435), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n491), .B2(new_n435), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n493), .A2(new_n494), .A3(new_n416), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n487), .B1(new_n495), .B2(new_n436), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n344), .A2(KEYINPUT85), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n341), .A2(new_n498), .A3(new_n343), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n493), .B2(new_n494), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n341), .A2(new_n343), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n461), .A2(new_n455), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(new_n452), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT39), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n476), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n467), .A2(new_n452), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT40), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n507), .B2(new_n509), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n511), .A2(new_n478), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n435), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n427), .A2(new_n429), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n421), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT38), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n427), .B2(new_n429), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n520), .B2(KEYINPUT86), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n421), .B1(new_n516), .B2(KEYINPUT37), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n523));
  AOI211_X1 g322(.A(new_n523), .B(new_n519), .C1(new_n427), .C2(new_n429), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n484), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT38), .B1(new_n522), .B2(new_n520), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n522), .A2(new_n524), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT87), .B1(new_n530), .B2(new_n521), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n414), .A2(new_n415), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT36), .ZN(new_n535));
  INV_X1    g334(.A(new_n415), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n536), .A2(KEYINPUT36), .A3(new_n413), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n501), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n284), .B1(new_n496), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n267), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n210), .B(new_n215), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT90), .B1(new_n545), .B2(new_n217), .ZN(new_n546));
  INV_X1    g345(.A(new_n222), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n212), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n267), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n262), .A2(new_n264), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n550), .B(new_n212), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  AOI211_X1 g350(.A(KEYINPUT97), .B(new_n544), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n268), .B2(new_n223), .ZN(new_n554));
  INV_X1    g353(.A(new_n544), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n543), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n543), .B(KEYINPUT99), .C1(new_n552), .C2(new_n556), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n560), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n549), .A2(new_n563), .A3(new_n551), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT100), .Z(new_n565));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n557), .A2(new_n560), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n565), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  INV_X1    g374(.A(new_n207), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n251), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n207), .A2(new_n250), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n207), .B(new_n250), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(KEYINPUT13), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n577), .A2(KEYINPUT18), .A3(new_n578), .A4(new_n580), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G197gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT11), .B(G169gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT88), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT12), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n582), .A3(new_n586), .A4(new_n587), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n574), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n540), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n491), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n203), .ZN(G1324gat));
  NOR2_X1   g402(.A1(new_n601), .A2(new_n435), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT42), .Z(new_n607));
  INV_X1    g406(.A(G8gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(new_n604), .ZN(G1325gat));
  INV_X1    g408(.A(G15gat), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n601), .A2(new_n610), .A3(new_n538), .ZN(new_n611));
  INV_X1    g410(.A(new_n534), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n540), .A2(new_n600), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n610), .B2(new_n613), .ZN(G1326gat));
  INV_X1    g413(.A(new_n500), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n601), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT43), .B(G22gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(G1327gat));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n496), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n491), .A2(new_n435), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT80), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n491), .A2(new_n492), .A3(new_n435), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n536), .A2(new_n413), .B1(new_n341), .B2(new_n343), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(KEYINPUT101), .A3(new_n487), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n539), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT44), .B1(new_n628), .B2(new_n282), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n239), .A2(new_n600), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n283), .B1(new_n496), .B2(new_n539), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(KEYINPUT44), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(G29gat), .B1(new_n634), .B2(new_n491), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G29gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n491), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT45), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n641), .ZN(G1328gat));
  OAI21_X1  g441(.A(G36gat), .B1(new_n634), .B2(new_n435), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n418), .A3(new_n514), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT46), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(G1329gat));
  INV_X1    g445(.A(new_n538), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n633), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n534), .A2(G43gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n648), .A2(G43gat), .B1(new_n637), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT101), .B1(new_n626), .B2(new_n487), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n619), .B(new_n486), .C1(new_n625), .C2(KEYINPUT35), .ZN(new_n654));
  INV_X1    g453(.A(new_n539), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n652), .B1(new_n656), .B2(new_n283), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n631), .A2(KEYINPUT44), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n657), .A2(new_n502), .A3(new_n636), .A4(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n628), .A2(new_n282), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n632), .B1(new_n662), .B2(new_n652), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n663), .A2(KEYINPUT104), .A3(new_n502), .A4(new_n636), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(G50gat), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT48), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n615), .A2(G50gat), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n637), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n665), .A2(new_n674), .ZN(new_n675));
  NOR4_X1   g474(.A1(new_n629), .A2(new_n632), .A3(new_n615), .A4(new_n630), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n670), .B1(new_n676), .B2(new_n336), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n666), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(KEYINPUT105), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1331gat));
  NOR2_X1   g482(.A1(new_n284), .A2(new_n598), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n628), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n574), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n639), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g488(.A(new_n435), .B(KEYINPUT107), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(KEYINPUT106), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n685), .A2(new_n693), .A3(new_n574), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  AND2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n687), .A2(new_n700), .A3(new_n612), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n538), .B1(new_n692), .B2(new_n694), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT50), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1334gat));
  AOI21_X1  g504(.A(new_n615), .B1(new_n692), .B2(new_n694), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g506(.A1(new_n240), .A2(new_n598), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n663), .A2(new_n574), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n253), .A3(new_n491), .ZN(new_n710));
  INV_X1    g509(.A(new_n662), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n708), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n708), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(KEYINPUT108), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n715), .A2(KEYINPUT108), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n639), .A4(new_n574), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n710), .B1(new_n718), .B2(new_n253), .ZN(G1336gat));
  INV_X1    g518(.A(new_n709), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n254), .B1(new_n720), .B2(new_n514), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n714), .A2(new_n715), .ZN(new_n722));
  INV_X1    g521(.A(new_n574), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n691), .A2(G92gat), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n691), .A2(G92gat), .ZN(new_n727));
  AND4_X1   g526(.A1(new_n574), .A2(new_n716), .A3(new_n717), .A4(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G92gat), .B1(new_n709), .B2(new_n691), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n726), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n725), .A2(new_n726), .B1(new_n728), .B2(new_n730), .ZN(G1337gat));
  NOR2_X1   g530(.A1(new_n534), .A2(G99gat), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n574), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G99gat), .B1(new_n709), .B2(new_n538), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1338gat));
  NOR3_X1   g537(.A1(new_n344), .A2(new_n723), .A3(G106gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n716), .A2(new_n717), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(G106gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n720), .B2(new_n502), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n720), .A2(new_n500), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n745), .A2(G106gat), .B1(new_n722), .B2(new_n739), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n742), .A2(new_n744), .B1(new_n746), .B2(new_n741), .ZN(G1339gat));
  OR2_X1    g546(.A1(new_n552), .A2(new_n556), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n749), .A3(new_n563), .A4(new_n543), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT110), .B1(new_n557), .B2(new_n560), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n562), .A2(KEYINPUT54), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n571), .A2(KEYINPUT54), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n569), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n752), .A2(KEYINPUT55), .A3(new_n754), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n570), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT55), .B1(new_n752), .B2(new_n754), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n759), .A2(new_n761), .A3(new_n598), .A4(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n579), .B2(new_n581), .ZN(new_n766));
  AOI211_X1 g565(.A(KEYINPUT112), .B(new_n580), .C1(new_n577), .C2(new_n578), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n583), .A2(new_n585), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n597), .B1(new_n769), .B2(new_n592), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n573), .B2(new_n570), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n282), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n759), .A2(new_n761), .A3(new_n282), .A4(new_n763), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n770), .B(KEYINPUT113), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n239), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NOR4_X1   g576(.A1(new_n239), .A2(new_n574), .A3(new_n598), .A4(new_n282), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n534), .B(new_n500), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n690), .A2(new_n491), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n376), .B1(new_n782), .B2(new_n598), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT114), .Z(new_n784));
  AOI21_X1  g583(.A(new_n491), .B1(new_n777), .B2(new_n779), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n624), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n690), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n376), .A3(new_n598), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n788), .ZN(G1340gat));
  INV_X1    g588(.A(new_n782), .ZN(new_n790));
  OAI21_X1  g589(.A(G120gat), .B1(new_n790), .B2(new_n723), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n574), .A2(new_n378), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT115), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n787), .B2(new_n240), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n240), .A2(G127gat), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n782), .B2(new_n797), .ZN(G1342gat));
  NOR4_X1   g597(.A1(new_n786), .A2(G134gat), .A3(new_n514), .A4(new_n283), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT116), .Z(new_n802));
  OAI21_X1  g601(.A(G134gat), .B1(new_n790), .B2(new_n283), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n802), .B(new_n803), .C1(new_n800), .C2(new_n799), .ZN(G1343gat));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n538), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n762), .A2(new_n599), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n771), .B1(new_n761), .B2(new_n808), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n774), .A2(new_n775), .B1(new_n809), .B2(new_n282), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n778), .B1(new_n810), .B2(new_n239), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n615), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT117), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n761), .A2(new_n808), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n283), .B1(new_n817), .B2(new_n771), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n762), .B(new_n758), .ZN(new_n819));
  INV_X1    g618(.A(new_n775), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n282), .A3(new_n761), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n240), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n816), .B(new_n813), .C1(new_n822), .C2(new_n778), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n777), .A2(new_n779), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n825), .B2(new_n502), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n598), .B(new_n807), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G141gat), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n647), .A2(new_n344), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n785), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT120), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n691), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n598), .A2(new_n305), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n805), .B(new_n828), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n830), .A2(new_n690), .A3(new_n833), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n827), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(KEYINPUT119), .A3(KEYINPUT58), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT119), .B1(new_n839), .B2(KEYINPUT58), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n834), .B1(new_n840), .B2(new_n841), .ZN(G1344gat));
  INV_X1    g641(.A(new_n832), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n307), .A3(new_n574), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n500), .B1(new_n811), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n822), .A2(KEYINPUT121), .A3(new_n778), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n812), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT122), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n825), .A2(KEYINPUT57), .A3(new_n502), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(KEYINPUT122), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n574), .A3(new_n807), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n845), .B1(new_n854), .B2(G148gat), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n824), .A2(new_n826), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n806), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT59), .B(new_n307), .C1(new_n857), .C2(new_n574), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n844), .B1(new_n855), .B2(new_n858), .ZN(G1345gat));
  AOI21_X1  g658(.A(G155gat), .B1(new_n843), .B2(new_n240), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n240), .A2(G155gat), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT123), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n857), .B2(new_n862), .ZN(G1346gat));
  NAND4_X1  g662(.A1(new_n831), .A2(new_n296), .A3(new_n435), .A4(new_n282), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n856), .A2(new_n283), .A3(new_n806), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n296), .B2(new_n865), .ZN(G1347gat));
  AOI211_X1 g665(.A(new_n639), .B(new_n691), .C1(new_n777), .C2(new_n779), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n624), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT124), .ZN(new_n869));
  INV_X1    g668(.A(G169gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n598), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n639), .A2(new_n435), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n780), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873), .B2(new_n599), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(G1348gat));
  INV_X1    g677(.A(G176gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n873), .A2(new_n879), .A3(new_n723), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n869), .A2(new_n574), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n879), .ZN(G1349gat));
  NAND3_X1  g681(.A1(new_n868), .A2(new_n350), .A3(new_n240), .ZN(new_n883));
  OAI21_X1  g682(.A(G183gat), .B1(new_n873), .B2(new_n239), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g684(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n351), .A3(new_n282), .ZN(new_n888));
  OAI21_X1  g687(.A(G190gat), .B1(new_n873), .B2(new_n283), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(KEYINPUT61), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(KEYINPUT61), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1351gat));
  XOR2_X1   g691(.A(KEYINPUT127), .B(G197gat), .Z(new_n893));
  AND2_X1   g692(.A1(new_n538), .A2(new_n872), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n853), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(new_n599), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n867), .A2(new_n829), .ZN(new_n897));
  INV_X1    g696(.A(new_n893), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n598), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1352gat));
  INV_X1    g699(.A(G204gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n901), .A3(new_n574), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT62), .Z(new_n903));
  AND3_X1   g702(.A1(new_n853), .A2(new_n574), .A3(new_n894), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n901), .ZN(G1353gat));
  NAND3_X1  g704(.A1(new_n897), .A2(new_n225), .A3(new_n240), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n853), .A2(new_n240), .A3(new_n894), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT63), .B1(new_n907), .B2(G211gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1354gat));
  OAI21_X1  g709(.A(G218gat), .B1(new_n895), .B2(new_n283), .ZN(new_n911));
  INV_X1    g710(.A(G218gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n912), .A3(new_n282), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1355gat));
endmodule


